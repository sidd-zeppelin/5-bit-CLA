magic
tech scmos
timestamp 1764717329
<< nwell >>
rect 58 69 90 101
rect 131 90 155 122
rect 209 69 241 101
rect 282 90 306 122
rect 58 4 110 36
rect 141 26 165 58
rect 220 4 272 36
rect 303 26 327 58
rect 466 57 498 89
rect 375 23 407 55
rect 466 1 498 33
rect 562 23 594 55
rect 58 -63 90 -31
rect 131 -42 155 -10
rect 200 -60 232 -20
rect 282 -42 306 -10
rect 330 -63 362 -31
rect 403 -42 427 -10
rect 457 -61 529 -21
rect 559 -42 583 -10
rect 720 -53 752 -21
rect 58 -128 110 -96
rect 141 -106 165 -74
rect 629 -87 661 -55
rect 58 -195 90 -163
rect 131 -174 155 -142
rect 210 -147 242 -99
rect 302 -124 326 -92
rect 350 -142 382 -102
rect 432 -124 456 -92
rect 476 -145 508 -113
rect 549 -124 573 -92
rect 720 -109 752 -77
rect 816 -87 848 -55
rect 597 -174 689 -126
rect 720 -153 744 -121
rect 873 -163 905 -131
rect 782 -197 814 -165
rect 58 -260 110 -228
rect 141 -238 165 -206
rect 213 -263 245 -207
rect 291 -231 315 -199
rect 343 -263 375 -215
rect 435 -240 459 -208
rect 483 -249 515 -209
rect 565 -231 589 -199
rect 615 -252 647 -220
rect 688 -231 712 -199
rect 873 -219 905 -187
rect 969 -197 1001 -165
rect 58 -327 90 -295
rect 131 -306 155 -274
rect 736 -292 848 -236
rect 877 -259 901 -227
rect 1034 -272 1066 -240
rect 943 -306 975 -274
rect 58 -392 110 -360
rect 141 -370 165 -338
rect 250 -383 273 -319
rect 332 -350 356 -318
rect 380 -371 412 -315
rect 458 -339 482 -307
rect 512 -362 544 -314
rect 604 -339 629 -307
rect 662 -357 694 -317
rect 744 -339 768 -307
rect 785 -360 817 -328
rect 858 -339 882 -307
rect 1034 -328 1066 -296
rect 1130 -306 1162 -274
rect 58 -460 90 -428
rect 131 -439 155 -407
rect 913 -413 1045 -349
rect 1083 -380 1107 -348
rect 1241 -383 1273 -351
rect 1150 -417 1182 -385
rect 1241 -439 1273 -407
rect 1337 -417 1369 -385
rect 58 -525 110 -493
rect 141 -503 165 -471
<< ntransistor >>
rect 97 88 117 90
rect 97 80 117 82
rect 248 88 268 90
rect 142 70 144 80
rect 248 80 268 82
rect 293 70 295 80
rect 508 76 528 78
rect 508 68 528 70
rect 417 42 437 44
rect 604 42 624 44
rect 417 34 437 36
rect 116 23 126 25
rect 116 15 126 17
rect 278 23 288 25
rect 152 6 154 16
rect 278 15 288 17
rect 604 34 624 36
rect 508 20 528 22
rect 314 6 316 16
rect 508 12 528 14
rect 238 -33 268 -31
rect 97 -44 117 -42
rect 97 -52 117 -50
rect 535 -34 545 -32
rect 238 -41 268 -39
rect 238 -49 268 -47
rect 142 -62 144 -52
rect 369 -44 389 -42
rect 293 -62 295 -52
rect 369 -52 389 -50
rect 762 -34 782 -32
rect 535 -42 545 -40
rect 535 -50 545 -48
rect 414 -62 416 -52
rect 762 -42 782 -40
rect 570 -62 572 -52
rect 671 -68 691 -66
rect 858 -68 878 -66
rect 671 -76 691 -74
rect 858 -76 878 -74
rect 762 -90 782 -88
rect 116 -109 126 -107
rect 116 -117 126 -115
rect 248 -112 288 -110
rect 152 -126 154 -116
rect 388 -115 418 -113
rect 248 -120 288 -118
rect 248 -128 288 -126
rect 248 -136 288 -134
rect 762 -98 782 -96
rect 388 -123 418 -121
rect 388 -131 418 -129
rect 313 -144 315 -134
rect 515 -126 535 -124
rect 443 -144 445 -134
rect 515 -134 535 -132
rect 560 -144 562 -134
rect 695 -139 705 -137
rect 695 -147 705 -145
rect 915 -144 935 -142
rect 695 -155 705 -153
rect 695 -163 705 -161
rect 915 -152 935 -150
rect 97 -176 117 -174
rect 97 -184 117 -182
rect 731 -173 733 -163
rect 824 -178 844 -176
rect 142 -194 144 -184
rect 1011 -178 1031 -176
rect 824 -186 844 -184
rect 1011 -186 1031 -184
rect 915 -200 935 -198
rect 251 -220 276 -218
rect 251 -228 276 -226
rect 116 -241 126 -239
rect 116 -249 126 -247
rect 251 -236 276 -234
rect 381 -228 421 -226
rect 521 -222 551 -220
rect 915 -208 935 -206
rect 521 -230 551 -228
rect 381 -236 421 -234
rect 251 -244 276 -242
rect 152 -258 154 -248
rect 251 -252 276 -250
rect 302 -251 304 -241
rect 381 -244 421 -242
rect 521 -238 551 -236
rect 654 -233 674 -231
rect 381 -252 421 -250
rect 446 -260 448 -250
rect 576 -251 578 -241
rect 654 -241 674 -239
rect 699 -251 701 -241
rect 854 -249 864 -247
rect 854 -257 864 -255
rect 854 -265 864 -263
rect 1076 -253 1096 -251
rect 1076 -261 1096 -259
rect 854 -273 864 -271
rect 888 -279 890 -269
rect 854 -281 864 -279
rect 985 -287 1005 -285
rect 1172 -287 1192 -285
rect 985 -295 1005 -293
rect 1172 -295 1192 -293
rect 97 -308 117 -306
rect 97 -316 117 -314
rect 1076 -309 1096 -307
rect 142 -326 144 -316
rect 281 -332 311 -330
rect 281 -340 311 -338
rect 418 -328 443 -326
rect 550 -327 590 -325
rect 418 -336 443 -334
rect 281 -348 311 -346
rect 281 -356 311 -354
rect 116 -373 126 -371
rect 116 -381 126 -379
rect 418 -344 443 -342
rect 700 -330 730 -328
rect 550 -335 590 -333
rect 550 -343 590 -341
rect 418 -352 443 -350
rect 281 -364 311 -362
rect 343 -370 345 -360
rect 418 -360 443 -358
rect 469 -359 471 -349
rect 1076 -317 1096 -315
rect 700 -338 730 -336
rect 700 -346 730 -344
rect 550 -351 590 -349
rect 616 -359 618 -349
rect 824 -341 844 -339
rect 755 -359 757 -349
rect 824 -349 844 -347
rect 869 -359 871 -349
rect 1051 -362 1061 -360
rect 281 -372 311 -370
rect 1051 -370 1061 -368
rect 1283 -364 1303 -362
rect 1283 -372 1303 -370
rect 1051 -378 1061 -376
rect 152 -390 154 -380
rect 1051 -386 1061 -384
rect 1051 -394 1061 -392
rect 1094 -400 1096 -390
rect 1192 -398 1212 -396
rect 1051 -402 1061 -400
rect 1379 -398 1399 -396
rect 1192 -406 1212 -404
rect 1379 -406 1399 -404
rect 1283 -420 1303 -418
rect 1283 -428 1303 -426
rect 97 -441 117 -439
rect 97 -449 117 -447
rect 142 -459 144 -449
rect 116 -506 126 -504
rect 116 -514 126 -512
rect 152 -523 154 -513
<< ptransistor >>
rect 142 96 144 116
rect 293 96 295 116
rect 64 88 84 90
rect 64 80 84 82
rect 215 88 235 90
rect 215 80 235 82
rect 472 76 492 78
rect 472 68 492 70
rect 152 32 154 52
rect 314 32 316 52
rect 381 42 401 44
rect 568 42 588 44
rect 381 34 401 36
rect 64 23 104 25
rect 64 15 104 17
rect 226 23 266 25
rect 226 15 266 17
rect 568 34 588 36
rect 472 20 492 22
rect 472 12 492 14
rect 142 -36 144 -16
rect 206 -33 226 -31
rect 64 -44 84 -42
rect 64 -52 84 -50
rect 293 -36 295 -16
rect 414 -36 416 -16
rect 463 -34 523 -32
rect 206 -41 226 -39
rect 206 -49 226 -47
rect 336 -44 356 -42
rect 336 -52 356 -50
rect 570 -36 572 -16
rect 726 -34 746 -32
rect 463 -42 523 -40
rect 463 -50 523 -48
rect 726 -42 746 -40
rect 635 -68 655 -66
rect 822 -68 842 -66
rect 635 -76 655 -74
rect 152 -100 154 -80
rect 822 -76 842 -74
rect 726 -90 746 -88
rect 64 -109 104 -107
rect 64 -117 104 -115
rect 216 -112 236 -110
rect 313 -118 315 -98
rect 356 -115 376 -113
rect 216 -120 236 -118
rect 216 -128 236 -126
rect 216 -136 236 -134
rect 443 -118 445 -98
rect 560 -118 562 -98
rect 726 -98 746 -96
rect 356 -123 376 -121
rect 356 -131 376 -129
rect 482 -126 502 -124
rect 482 -134 502 -132
rect 603 -139 683 -137
rect 603 -147 683 -145
rect 731 -147 733 -127
rect 879 -144 899 -142
rect 142 -168 144 -148
rect 603 -155 683 -153
rect 603 -163 683 -161
rect 879 -152 899 -150
rect 64 -176 84 -174
rect 64 -184 84 -182
rect 788 -178 808 -176
rect 975 -178 995 -176
rect 788 -186 808 -184
rect 975 -186 995 -184
rect 879 -200 899 -198
rect 152 -232 154 -212
rect 219 -220 239 -218
rect 302 -225 304 -205
rect 219 -228 239 -226
rect 64 -241 104 -239
rect 64 -249 104 -247
rect 219 -236 239 -234
rect 349 -228 369 -226
rect 446 -234 448 -214
rect 489 -222 509 -220
rect 576 -225 578 -205
rect 699 -225 701 -205
rect 879 -208 899 -206
rect 489 -230 509 -228
rect 349 -236 369 -234
rect 219 -244 239 -242
rect 219 -252 239 -250
rect 349 -244 369 -242
rect 489 -238 509 -236
rect 621 -233 641 -231
rect 349 -252 369 -250
rect 621 -241 641 -239
rect 742 -249 842 -247
rect 888 -253 890 -233
rect 742 -257 842 -255
rect 742 -265 842 -263
rect 1040 -253 1060 -251
rect 1040 -261 1060 -259
rect 742 -273 842 -271
rect 142 -300 144 -280
rect 742 -281 842 -279
rect 949 -287 969 -285
rect 1136 -287 1156 -285
rect 949 -295 969 -293
rect 1136 -295 1156 -293
rect 64 -308 84 -306
rect 64 -316 84 -314
rect 1040 -309 1060 -307
rect 257 -332 267 -330
rect 257 -340 267 -338
rect 152 -364 154 -344
rect 343 -344 345 -324
rect 386 -328 406 -326
rect 469 -333 471 -313
rect 518 -327 538 -325
rect 386 -336 406 -334
rect 257 -348 267 -346
rect 257 -356 267 -354
rect 64 -373 104 -371
rect 64 -381 104 -379
rect 386 -344 406 -342
rect 616 -333 618 -313
rect 668 -330 688 -328
rect 518 -335 538 -333
rect 518 -343 538 -341
rect 386 -352 406 -350
rect 257 -364 267 -362
rect 386 -360 406 -358
rect 755 -333 757 -313
rect 869 -333 871 -313
rect 1040 -317 1060 -315
rect 668 -338 688 -336
rect 668 -346 688 -344
rect 518 -351 538 -349
rect 791 -341 811 -339
rect 791 -349 811 -347
rect 919 -362 1039 -360
rect 257 -372 267 -370
rect 919 -370 1039 -368
rect 1094 -374 1096 -354
rect 1247 -364 1267 -362
rect 1247 -372 1267 -370
rect 919 -378 1039 -376
rect 919 -386 1039 -384
rect 919 -394 1039 -392
rect 1156 -398 1176 -396
rect 919 -402 1039 -400
rect 1343 -398 1363 -396
rect 1156 -406 1176 -404
rect 1343 -406 1363 -404
rect 142 -433 144 -413
rect 1247 -420 1267 -418
rect 1247 -428 1267 -426
rect 64 -441 84 -439
rect 64 -449 84 -447
rect 152 -497 154 -477
rect 64 -506 104 -504
rect 64 -514 104 -512
<< ndiffusion >>
rect 97 90 117 91
rect 97 87 117 88
rect 97 82 117 83
rect 248 90 268 91
rect 97 79 117 80
rect 141 70 142 80
rect 144 70 145 80
rect 248 87 268 88
rect 248 82 268 83
rect 248 79 268 80
rect 292 70 293 80
rect 295 70 296 80
rect 508 78 528 79
rect 508 75 528 76
rect 508 70 528 71
rect 508 67 528 68
rect 417 44 437 45
rect 417 41 437 42
rect 604 44 624 45
rect 417 36 437 37
rect 116 25 126 26
rect 116 22 126 23
rect 116 17 126 18
rect 278 25 288 26
rect 116 14 126 15
rect 151 6 152 16
rect 154 6 155 16
rect 278 22 288 23
rect 278 17 288 18
rect 417 33 437 34
rect 604 41 624 42
rect 604 36 624 37
rect 604 33 624 34
rect 508 22 528 23
rect 278 14 288 15
rect 313 6 314 16
rect 316 6 317 16
rect 508 19 528 20
rect 508 14 528 15
rect 508 11 528 12
rect 238 -31 268 -30
rect 97 -42 117 -41
rect 97 -45 117 -44
rect 97 -50 117 -49
rect 238 -34 268 -33
rect 535 -32 545 -31
rect 238 -39 268 -38
rect 238 -42 268 -41
rect 238 -47 268 -46
rect 97 -53 117 -52
rect 141 -62 142 -52
rect 144 -62 145 -52
rect 238 -50 268 -49
rect 369 -42 389 -41
rect 292 -62 293 -52
rect 295 -62 296 -52
rect 369 -45 389 -44
rect 369 -50 389 -49
rect 535 -35 545 -34
rect 762 -32 782 -31
rect 535 -40 545 -39
rect 535 -43 545 -42
rect 535 -48 545 -47
rect 369 -53 389 -52
rect 413 -62 414 -52
rect 416 -62 417 -52
rect 535 -51 545 -50
rect 762 -35 782 -34
rect 762 -40 782 -39
rect 762 -43 782 -42
rect 569 -62 570 -52
rect 572 -62 573 -52
rect 671 -66 691 -65
rect 671 -69 691 -68
rect 858 -66 878 -65
rect 671 -74 691 -73
rect 671 -77 691 -76
rect 858 -69 878 -68
rect 858 -74 878 -73
rect 858 -77 878 -76
rect 762 -88 782 -87
rect 116 -107 126 -106
rect 116 -110 126 -109
rect 116 -115 126 -114
rect 248 -110 288 -109
rect 116 -118 126 -117
rect 151 -126 152 -116
rect 154 -126 155 -116
rect 248 -113 288 -112
rect 248 -118 288 -117
rect 388 -113 418 -112
rect 248 -121 288 -120
rect 248 -126 288 -125
rect 248 -129 288 -128
rect 248 -134 288 -133
rect 248 -137 288 -136
rect 388 -116 418 -115
rect 762 -91 782 -90
rect 762 -96 782 -95
rect 762 -99 782 -98
rect 388 -121 418 -120
rect 388 -124 418 -123
rect 388 -129 418 -128
rect 312 -144 313 -134
rect 315 -144 316 -134
rect 388 -132 418 -131
rect 515 -124 535 -123
rect 442 -144 443 -134
rect 445 -144 446 -134
rect 515 -127 535 -126
rect 515 -132 535 -131
rect 515 -135 535 -134
rect 559 -144 560 -134
rect 562 -144 563 -134
rect 695 -137 705 -136
rect 695 -140 705 -139
rect 695 -145 705 -144
rect 915 -142 935 -141
rect 695 -148 705 -147
rect 695 -153 705 -152
rect 695 -156 705 -155
rect 695 -161 705 -160
rect 915 -145 935 -144
rect 915 -150 935 -149
rect 915 -153 935 -152
rect 695 -164 705 -163
rect 97 -174 117 -173
rect 97 -177 117 -176
rect 97 -182 117 -181
rect 730 -173 731 -163
rect 733 -173 734 -163
rect 824 -176 844 -175
rect 97 -185 117 -184
rect 141 -194 142 -184
rect 144 -194 145 -184
rect 824 -179 844 -178
rect 1011 -176 1031 -175
rect 824 -184 844 -183
rect 824 -187 844 -186
rect 1011 -179 1031 -178
rect 1011 -184 1031 -183
rect 1011 -187 1031 -186
rect 915 -198 935 -197
rect 251 -218 276 -217
rect 251 -221 276 -220
rect 251 -226 276 -225
rect 116 -239 126 -238
rect 116 -242 126 -241
rect 116 -247 126 -246
rect 251 -229 276 -228
rect 251 -234 276 -233
rect 251 -237 276 -236
rect 381 -226 421 -225
rect 381 -229 421 -228
rect 381 -234 421 -233
rect 521 -220 551 -219
rect 521 -223 551 -222
rect 915 -201 935 -200
rect 915 -206 935 -205
rect 915 -209 935 -208
rect 521 -228 551 -227
rect 251 -242 276 -241
rect 116 -250 126 -249
rect 151 -258 152 -248
rect 154 -258 155 -248
rect 251 -245 276 -244
rect 251 -250 276 -249
rect 301 -251 302 -241
rect 304 -251 305 -241
rect 381 -237 421 -236
rect 381 -242 421 -241
rect 251 -253 276 -252
rect 381 -245 421 -244
rect 381 -250 421 -249
rect 521 -231 551 -230
rect 521 -236 551 -235
rect 521 -239 551 -238
rect 654 -231 674 -230
rect 381 -253 421 -252
rect 445 -260 446 -250
rect 448 -260 449 -250
rect 575 -251 576 -241
rect 578 -251 579 -241
rect 654 -234 674 -233
rect 654 -239 674 -238
rect 654 -242 674 -241
rect 698 -251 699 -241
rect 701 -251 702 -241
rect 854 -247 864 -246
rect 854 -250 864 -249
rect 854 -255 864 -254
rect 854 -258 864 -257
rect 854 -263 864 -262
rect 854 -266 864 -265
rect 1076 -251 1096 -250
rect 1076 -254 1096 -253
rect 1076 -259 1096 -258
rect 1076 -262 1096 -261
rect 854 -271 864 -270
rect 854 -274 864 -273
rect 854 -279 864 -278
rect 887 -279 888 -269
rect 890 -279 891 -269
rect 854 -282 864 -281
rect 985 -285 1005 -284
rect 985 -288 1005 -287
rect 1172 -285 1192 -284
rect 985 -293 1005 -292
rect 985 -296 1005 -295
rect 1172 -288 1192 -287
rect 1172 -293 1192 -292
rect 1172 -296 1192 -295
rect 97 -306 117 -305
rect 97 -309 117 -308
rect 97 -314 117 -313
rect 1076 -307 1096 -306
rect 97 -317 117 -316
rect 141 -326 142 -316
rect 144 -326 145 -316
rect 281 -330 311 -329
rect 281 -333 311 -332
rect 281 -338 311 -337
rect 281 -341 311 -340
rect 418 -326 443 -325
rect 418 -329 443 -328
rect 550 -325 590 -324
rect 418 -334 443 -333
rect 281 -346 311 -345
rect 281 -349 311 -348
rect 281 -354 311 -353
rect 116 -371 126 -370
rect 116 -374 126 -373
rect 116 -379 126 -378
rect 281 -357 311 -356
rect 418 -337 443 -336
rect 418 -342 443 -341
rect 418 -345 443 -344
rect 550 -328 590 -327
rect 550 -333 590 -332
rect 700 -328 730 -327
rect 550 -336 590 -335
rect 550 -341 590 -340
rect 418 -350 443 -349
rect 281 -362 311 -361
rect 281 -365 311 -364
rect 281 -370 311 -369
rect 342 -370 343 -360
rect 345 -370 346 -360
rect 418 -353 443 -352
rect 418 -358 443 -357
rect 468 -359 469 -349
rect 471 -359 472 -349
rect 550 -344 590 -343
rect 550 -349 590 -348
rect 700 -331 730 -330
rect 1076 -310 1096 -309
rect 1076 -315 1096 -314
rect 1076 -318 1096 -317
rect 700 -336 730 -335
rect 700 -339 730 -338
rect 700 -344 730 -343
rect 550 -352 590 -351
rect 615 -359 616 -349
rect 618 -359 619 -349
rect 700 -347 730 -346
rect 824 -339 844 -338
rect 754 -359 755 -349
rect 757 -359 758 -349
rect 824 -342 844 -341
rect 824 -347 844 -346
rect 824 -350 844 -349
rect 868 -359 869 -349
rect 871 -359 872 -349
rect 418 -361 443 -360
rect 1051 -360 1061 -359
rect 281 -373 311 -372
rect 1051 -363 1061 -362
rect 1051 -368 1061 -367
rect 1051 -371 1061 -370
rect 1283 -362 1303 -361
rect 1283 -365 1303 -364
rect 1283 -370 1303 -369
rect 1051 -376 1061 -375
rect 116 -382 126 -381
rect 151 -390 152 -380
rect 154 -390 155 -380
rect 1051 -379 1061 -378
rect 1051 -384 1061 -383
rect 1051 -387 1061 -386
rect 1283 -373 1303 -372
rect 1051 -392 1061 -391
rect 1051 -395 1061 -394
rect 1051 -400 1061 -399
rect 1093 -400 1094 -390
rect 1096 -400 1097 -390
rect 1192 -396 1212 -395
rect 1051 -403 1061 -402
rect 1192 -399 1212 -398
rect 1379 -396 1399 -395
rect 1192 -404 1212 -403
rect 1192 -407 1212 -406
rect 1379 -399 1399 -398
rect 1379 -404 1399 -403
rect 1379 -407 1399 -406
rect 1283 -418 1303 -417
rect 1283 -421 1303 -420
rect 1283 -426 1303 -425
rect 1283 -429 1303 -428
rect 97 -439 117 -438
rect 97 -442 117 -441
rect 97 -447 117 -446
rect 97 -450 117 -449
rect 141 -459 142 -449
rect 144 -459 145 -449
rect 116 -504 126 -503
rect 116 -507 126 -506
rect 116 -512 126 -511
rect 116 -515 126 -514
rect 151 -523 152 -513
rect 154 -523 155 -513
<< pdiffusion >>
rect 141 96 142 116
rect 144 96 145 116
rect 292 96 293 116
rect 295 96 296 116
rect 64 90 84 91
rect 64 87 84 88
rect 64 82 84 83
rect 215 90 235 91
rect 215 87 235 88
rect 64 79 84 80
rect 215 82 235 83
rect 215 79 235 80
rect 472 78 492 79
rect 472 75 492 76
rect 472 70 492 71
rect 472 67 492 68
rect 151 32 152 52
rect 154 32 155 52
rect 313 32 314 52
rect 316 32 317 52
rect 381 44 401 45
rect 381 41 401 42
rect 381 36 401 37
rect 568 44 588 45
rect 568 41 588 42
rect 381 33 401 34
rect 64 25 104 26
rect 64 22 104 23
rect 64 17 104 18
rect 226 25 266 26
rect 226 22 266 23
rect 64 14 104 15
rect 226 17 266 18
rect 568 36 588 37
rect 568 33 588 34
rect 472 22 492 23
rect 472 19 492 20
rect 226 14 266 15
rect 472 14 492 15
rect 472 11 492 12
rect 141 -36 142 -16
rect 144 -36 145 -16
rect 206 -31 226 -30
rect 206 -34 226 -33
rect 64 -42 84 -41
rect 64 -45 84 -44
rect 64 -50 84 -49
rect 206 -39 226 -38
rect 292 -36 293 -16
rect 295 -36 296 -16
rect 413 -36 414 -16
rect 416 -36 417 -16
rect 463 -32 523 -31
rect 463 -35 523 -34
rect 206 -42 226 -41
rect 206 -47 226 -46
rect 206 -50 226 -49
rect 64 -53 84 -52
rect 336 -42 356 -41
rect 336 -45 356 -44
rect 336 -50 356 -49
rect 463 -40 523 -39
rect 569 -36 570 -16
rect 572 -36 573 -16
rect 726 -32 746 -31
rect 726 -35 746 -34
rect 463 -43 523 -42
rect 463 -48 523 -47
rect 463 -51 523 -50
rect 336 -53 356 -52
rect 726 -40 746 -39
rect 726 -43 746 -42
rect 635 -66 655 -65
rect 635 -69 655 -68
rect 635 -74 655 -73
rect 822 -66 842 -65
rect 822 -69 842 -68
rect 635 -77 655 -76
rect 151 -100 152 -80
rect 154 -100 155 -80
rect 822 -74 842 -73
rect 822 -77 842 -76
rect 726 -88 746 -87
rect 726 -91 746 -90
rect 64 -107 104 -106
rect 64 -110 104 -109
rect 64 -115 104 -114
rect 216 -110 236 -109
rect 216 -113 236 -112
rect 64 -118 104 -117
rect 216 -118 236 -117
rect 312 -118 313 -98
rect 315 -118 316 -98
rect 356 -113 376 -112
rect 356 -116 376 -115
rect 216 -121 236 -120
rect 216 -126 236 -125
rect 216 -129 236 -128
rect 216 -134 236 -133
rect 216 -137 236 -136
rect 356 -121 376 -120
rect 442 -118 443 -98
rect 445 -118 446 -98
rect 559 -118 560 -98
rect 562 -118 563 -98
rect 726 -96 746 -95
rect 726 -99 746 -98
rect 356 -124 376 -123
rect 356 -129 376 -128
rect 356 -132 376 -131
rect 482 -124 502 -123
rect 482 -127 502 -126
rect 482 -132 502 -131
rect 482 -135 502 -134
rect 603 -137 683 -136
rect 603 -140 683 -139
rect 603 -145 683 -144
rect 730 -147 731 -127
rect 733 -147 734 -127
rect 879 -142 899 -141
rect 879 -145 899 -144
rect 603 -148 683 -147
rect 141 -168 142 -148
rect 144 -168 145 -148
rect 603 -153 683 -152
rect 603 -156 683 -155
rect 603 -161 683 -160
rect 879 -150 899 -149
rect 879 -153 899 -152
rect 603 -164 683 -163
rect 64 -174 84 -173
rect 64 -177 84 -176
rect 64 -182 84 -181
rect 788 -176 808 -175
rect 788 -179 808 -178
rect 64 -185 84 -184
rect 788 -184 808 -183
rect 975 -176 995 -175
rect 975 -179 995 -178
rect 788 -187 808 -186
rect 975 -184 995 -183
rect 975 -187 995 -186
rect 879 -198 899 -197
rect 879 -201 899 -200
rect 151 -232 152 -212
rect 154 -232 155 -212
rect 219 -218 239 -217
rect 219 -221 239 -220
rect 219 -226 239 -225
rect 301 -225 302 -205
rect 304 -225 305 -205
rect 219 -229 239 -228
rect 64 -239 104 -238
rect 64 -242 104 -241
rect 64 -247 104 -246
rect 219 -234 239 -233
rect 219 -237 239 -236
rect 219 -242 239 -241
rect 349 -226 369 -225
rect 349 -229 369 -228
rect 349 -234 369 -233
rect 445 -234 446 -214
rect 448 -234 449 -214
rect 489 -220 509 -219
rect 489 -223 509 -222
rect 489 -228 509 -227
rect 575 -225 576 -205
rect 578 -225 579 -205
rect 698 -225 699 -205
rect 701 -225 702 -205
rect 879 -206 899 -205
rect 879 -209 899 -208
rect 489 -231 509 -230
rect 349 -237 369 -236
rect 219 -245 239 -244
rect 64 -250 104 -249
rect 219 -250 239 -249
rect 349 -242 369 -241
rect 349 -245 369 -244
rect 219 -253 239 -252
rect 349 -250 369 -249
rect 489 -236 509 -235
rect 489 -239 509 -238
rect 621 -231 641 -230
rect 621 -234 641 -233
rect 349 -253 369 -252
rect 621 -239 641 -238
rect 621 -242 641 -241
rect 742 -247 842 -246
rect 742 -250 842 -249
rect 742 -255 842 -254
rect 887 -253 888 -233
rect 890 -253 891 -233
rect 742 -258 842 -257
rect 742 -263 842 -262
rect 742 -266 842 -265
rect 742 -271 842 -270
rect 1040 -251 1060 -250
rect 1040 -254 1060 -253
rect 1040 -259 1060 -258
rect 1040 -262 1060 -261
rect 742 -274 842 -273
rect 141 -300 142 -280
rect 144 -300 145 -280
rect 742 -279 842 -278
rect 742 -282 842 -281
rect 949 -285 969 -284
rect 949 -288 969 -287
rect 949 -293 969 -292
rect 1136 -285 1156 -284
rect 1136 -288 1156 -287
rect 949 -296 969 -295
rect 1136 -293 1156 -292
rect 1136 -296 1156 -295
rect 64 -306 84 -305
rect 64 -309 84 -308
rect 64 -314 84 -313
rect 1040 -307 1060 -306
rect 1040 -310 1060 -309
rect 64 -317 84 -316
rect 257 -330 267 -329
rect 257 -333 267 -332
rect 257 -338 267 -337
rect 257 -341 267 -340
rect 151 -364 152 -344
rect 154 -364 155 -344
rect 257 -346 267 -345
rect 342 -344 343 -324
rect 345 -344 346 -324
rect 386 -326 406 -325
rect 386 -329 406 -328
rect 386 -334 406 -333
rect 468 -333 469 -313
rect 471 -333 472 -313
rect 518 -325 538 -324
rect 518 -328 538 -327
rect 386 -337 406 -336
rect 257 -349 267 -348
rect 257 -354 267 -353
rect 257 -357 267 -356
rect 64 -371 104 -370
rect 64 -374 104 -373
rect 64 -379 104 -378
rect 257 -362 267 -361
rect 386 -342 406 -341
rect 386 -345 406 -344
rect 386 -350 406 -349
rect 518 -333 538 -332
rect 615 -333 616 -313
rect 618 -333 619 -313
rect 668 -328 688 -327
rect 668 -331 688 -330
rect 518 -336 538 -335
rect 518 -341 538 -340
rect 518 -344 538 -343
rect 386 -353 406 -352
rect 257 -365 267 -364
rect 257 -370 267 -369
rect 386 -358 406 -357
rect 518 -349 538 -348
rect 668 -336 688 -335
rect 754 -333 755 -313
rect 757 -333 758 -313
rect 868 -333 869 -313
rect 871 -333 872 -313
rect 1040 -315 1060 -314
rect 1040 -318 1060 -317
rect 668 -339 688 -338
rect 668 -344 688 -343
rect 668 -347 688 -346
rect 518 -352 538 -351
rect 791 -339 811 -338
rect 791 -342 811 -341
rect 791 -347 811 -346
rect 791 -350 811 -349
rect 386 -361 406 -360
rect 919 -360 1039 -359
rect 919 -363 1039 -362
rect 257 -373 267 -372
rect 919 -368 1039 -367
rect 919 -371 1039 -370
rect 919 -376 1039 -375
rect 1093 -374 1094 -354
rect 1096 -374 1097 -354
rect 1247 -362 1267 -361
rect 1247 -365 1267 -364
rect 1247 -370 1267 -369
rect 1247 -373 1267 -372
rect 919 -379 1039 -378
rect 64 -382 104 -381
rect 919 -384 1039 -383
rect 919 -387 1039 -386
rect 919 -392 1039 -391
rect 919 -395 1039 -394
rect 919 -400 1039 -399
rect 1156 -396 1176 -395
rect 1156 -399 1176 -398
rect 919 -403 1039 -402
rect 1156 -404 1176 -403
rect 1343 -396 1363 -395
rect 1343 -399 1363 -398
rect 1156 -407 1176 -406
rect 1343 -404 1363 -403
rect 1343 -407 1363 -406
rect 141 -433 142 -413
rect 144 -433 145 -413
rect 1247 -418 1267 -417
rect 1247 -421 1267 -420
rect 1247 -426 1267 -425
rect 1247 -429 1267 -428
rect 64 -439 84 -438
rect 64 -442 84 -441
rect 64 -447 84 -446
rect 64 -450 84 -449
rect 151 -497 152 -477
rect 154 -497 155 -477
rect 64 -504 104 -503
rect 64 -507 104 -506
rect 64 -512 104 -511
rect 64 -515 104 -514
<< ndcontact >>
rect 97 91 117 95
rect 97 83 117 87
rect 248 91 268 95
rect 97 75 117 79
rect 137 70 141 80
rect 145 70 149 80
rect 248 83 268 87
rect 248 75 268 79
rect 288 70 292 80
rect 296 70 300 80
rect 508 79 528 83
rect 508 71 528 75
rect 508 63 528 67
rect 417 45 437 49
rect 604 45 624 49
rect 417 37 437 41
rect 116 26 126 30
rect 116 18 126 22
rect 278 26 288 30
rect 116 10 126 14
rect 147 6 151 16
rect 155 6 159 16
rect 278 18 288 22
rect 604 37 624 41
rect 417 29 437 33
rect 604 29 624 33
rect 508 23 528 27
rect 278 10 288 14
rect 309 6 313 16
rect 317 6 321 16
rect 508 15 528 19
rect 508 7 528 11
rect 238 -30 268 -26
rect 97 -41 117 -37
rect 97 -49 117 -45
rect 238 -38 268 -34
rect 535 -31 545 -27
rect 238 -46 268 -42
rect 97 -57 117 -53
rect 137 -62 141 -52
rect 145 -62 149 -52
rect 238 -54 268 -50
rect 369 -41 389 -37
rect 288 -62 292 -52
rect 296 -62 300 -52
rect 369 -49 389 -45
rect 535 -39 545 -35
rect 762 -31 782 -27
rect 535 -47 545 -43
rect 369 -57 389 -53
rect 409 -62 413 -52
rect 417 -62 421 -52
rect 535 -55 545 -51
rect 762 -39 782 -35
rect 762 -47 782 -43
rect 565 -62 569 -52
rect 573 -62 577 -52
rect 671 -65 691 -61
rect 858 -65 878 -61
rect 671 -73 691 -69
rect 858 -73 878 -69
rect 671 -81 691 -77
rect 858 -81 878 -77
rect 762 -87 782 -83
rect 116 -106 126 -102
rect 116 -114 126 -110
rect 248 -109 288 -105
rect 116 -122 126 -118
rect 147 -126 151 -116
rect 155 -126 159 -116
rect 248 -117 288 -113
rect 388 -112 418 -108
rect 248 -125 288 -121
rect 248 -133 288 -129
rect 248 -141 288 -137
rect 388 -120 418 -116
rect 762 -95 782 -91
rect 762 -103 782 -99
rect 388 -128 418 -124
rect 308 -144 312 -134
rect 316 -144 320 -134
rect 388 -136 418 -132
rect 515 -123 535 -119
rect 438 -144 442 -134
rect 446 -144 450 -134
rect 515 -131 535 -127
rect 515 -139 535 -135
rect 555 -144 559 -134
rect 563 -144 567 -134
rect 695 -136 705 -132
rect 695 -144 705 -140
rect 915 -141 935 -137
rect 695 -152 705 -148
rect 695 -160 705 -156
rect 915 -149 935 -145
rect 915 -157 935 -153
rect 695 -168 705 -164
rect 97 -173 117 -169
rect 97 -181 117 -177
rect 726 -173 730 -163
rect 734 -173 738 -163
rect 824 -175 844 -171
rect 97 -189 117 -185
rect 137 -194 141 -184
rect 145 -194 149 -184
rect 1011 -175 1031 -171
rect 824 -183 844 -179
rect 1011 -183 1031 -179
rect 824 -191 844 -187
rect 1011 -191 1031 -187
rect 915 -197 935 -193
rect 251 -217 276 -213
rect 251 -225 276 -221
rect 116 -238 126 -234
rect 116 -246 126 -242
rect 251 -233 276 -229
rect 251 -241 276 -237
rect 381 -225 421 -221
rect 381 -233 421 -229
rect 521 -219 551 -215
rect 521 -227 551 -223
rect 915 -205 935 -201
rect 915 -213 935 -209
rect 116 -254 126 -250
rect 147 -258 151 -248
rect 155 -258 159 -248
rect 251 -249 276 -245
rect 297 -251 301 -241
rect 305 -251 309 -241
rect 381 -241 421 -237
rect 251 -257 276 -253
rect 381 -249 421 -245
rect 521 -235 551 -231
rect 521 -243 551 -239
rect 654 -230 674 -226
rect 381 -257 421 -253
rect 441 -260 445 -250
rect 449 -260 453 -250
rect 571 -251 575 -241
rect 579 -251 583 -241
rect 654 -238 674 -234
rect 654 -246 674 -242
rect 694 -251 698 -241
rect 702 -251 706 -241
rect 854 -246 864 -242
rect 854 -254 864 -250
rect 854 -262 864 -258
rect 854 -270 864 -266
rect 1076 -250 1096 -246
rect 1076 -258 1096 -254
rect 1076 -266 1096 -262
rect 854 -278 864 -274
rect 883 -279 887 -269
rect 891 -279 895 -269
rect 854 -286 864 -282
rect 985 -284 1005 -280
rect 1172 -284 1192 -280
rect 985 -292 1005 -288
rect 1172 -292 1192 -288
rect 985 -300 1005 -296
rect 1172 -300 1192 -296
rect 97 -305 117 -301
rect 97 -313 117 -309
rect 1076 -306 1096 -302
rect 97 -321 117 -317
rect 137 -326 141 -316
rect 145 -326 149 -316
rect 281 -329 311 -325
rect 281 -337 311 -333
rect 281 -345 311 -341
rect 418 -325 443 -321
rect 418 -333 443 -329
rect 550 -324 590 -320
rect 281 -353 311 -349
rect 116 -370 126 -366
rect 116 -378 126 -374
rect 281 -361 311 -357
rect 418 -341 443 -337
rect 418 -349 443 -345
rect 550 -332 590 -328
rect 700 -327 730 -323
rect 550 -340 590 -336
rect 281 -369 311 -365
rect 338 -370 342 -360
rect 346 -370 350 -360
rect 418 -357 443 -353
rect 464 -359 468 -349
rect 472 -359 476 -349
rect 550 -348 590 -344
rect 700 -335 730 -331
rect 1076 -314 1096 -310
rect 1076 -322 1096 -318
rect 700 -343 730 -339
rect 550 -356 590 -352
rect 611 -359 615 -349
rect 619 -359 623 -349
rect 700 -351 730 -347
rect 824 -338 844 -334
rect 750 -359 754 -349
rect 758 -359 762 -349
rect 824 -346 844 -342
rect 824 -354 844 -350
rect 864 -359 868 -349
rect 872 -359 876 -349
rect 418 -365 443 -361
rect 1051 -359 1061 -355
rect 1051 -367 1061 -363
rect 281 -377 311 -373
rect 1051 -375 1061 -371
rect 1283 -361 1303 -357
rect 1283 -369 1303 -365
rect 116 -386 126 -382
rect 147 -390 151 -380
rect 155 -390 159 -380
rect 1051 -383 1061 -379
rect 1051 -391 1061 -387
rect 1283 -377 1303 -373
rect 1051 -399 1061 -395
rect 1089 -400 1093 -390
rect 1097 -400 1101 -390
rect 1192 -395 1212 -391
rect 1051 -407 1061 -403
rect 1379 -395 1399 -391
rect 1192 -403 1212 -399
rect 1379 -403 1399 -399
rect 1192 -411 1212 -407
rect 1379 -411 1399 -407
rect 1283 -417 1303 -413
rect 1283 -425 1303 -421
rect 1283 -433 1303 -429
rect 97 -438 117 -434
rect 97 -446 117 -442
rect 97 -454 117 -450
rect 137 -459 141 -449
rect 145 -459 149 -449
rect 116 -503 126 -499
rect 116 -511 126 -507
rect 116 -519 126 -515
rect 147 -523 151 -513
rect 155 -523 159 -513
<< pdcontact >>
rect 137 96 141 116
rect 145 96 149 116
rect 288 96 292 116
rect 296 96 300 116
rect 64 91 84 95
rect 64 83 84 87
rect 215 91 235 95
rect 215 83 235 87
rect 64 75 84 79
rect 215 75 235 79
rect 472 79 492 83
rect 472 71 492 75
rect 472 63 492 67
rect 147 32 151 52
rect 155 32 159 52
rect 309 32 313 52
rect 317 32 321 52
rect 381 45 401 49
rect 568 45 588 49
rect 381 37 401 41
rect 568 37 588 41
rect 64 26 104 30
rect 64 18 104 22
rect 226 26 266 30
rect 226 18 266 22
rect 64 10 104 14
rect 381 29 401 33
rect 568 29 588 33
rect 472 23 492 27
rect 226 10 266 14
rect 472 15 492 19
rect 472 7 492 11
rect 137 -36 141 -16
rect 145 -36 149 -16
rect 206 -30 226 -26
rect 64 -41 84 -37
rect 64 -49 84 -45
rect 206 -38 226 -34
rect 288 -36 292 -16
rect 296 -36 300 -16
rect 409 -36 413 -16
rect 417 -36 421 -16
rect 463 -31 523 -27
rect 206 -46 226 -42
rect 64 -57 84 -53
rect 206 -54 226 -50
rect 336 -41 356 -37
rect 336 -49 356 -45
rect 463 -39 523 -35
rect 565 -36 569 -16
rect 573 -36 577 -16
rect 726 -31 746 -27
rect 463 -47 523 -43
rect 336 -57 356 -53
rect 463 -55 523 -51
rect 726 -39 746 -35
rect 726 -47 746 -43
rect 635 -65 655 -61
rect 822 -65 842 -61
rect 635 -73 655 -69
rect 822 -73 842 -69
rect 147 -100 151 -80
rect 155 -100 159 -80
rect 635 -81 655 -77
rect 822 -81 842 -77
rect 726 -87 746 -83
rect 726 -95 746 -91
rect 64 -106 104 -102
rect 64 -114 104 -110
rect 216 -109 236 -105
rect 64 -122 104 -118
rect 216 -117 236 -113
rect 308 -118 312 -98
rect 316 -118 320 -98
rect 356 -112 376 -108
rect 216 -125 236 -121
rect 216 -133 236 -129
rect 216 -141 236 -137
rect 356 -120 376 -116
rect 438 -118 442 -98
rect 446 -118 450 -98
rect 555 -118 559 -98
rect 563 -118 567 -98
rect 726 -103 746 -99
rect 356 -128 376 -124
rect 356 -136 376 -132
rect 482 -123 502 -119
rect 482 -131 502 -127
rect 482 -139 502 -135
rect 603 -136 683 -132
rect 603 -144 683 -140
rect 726 -147 730 -127
rect 734 -147 738 -127
rect 879 -141 899 -137
rect 137 -168 141 -148
rect 145 -168 149 -148
rect 603 -152 683 -148
rect 603 -160 683 -156
rect 879 -149 899 -145
rect 879 -157 899 -153
rect 603 -168 683 -164
rect 64 -173 84 -169
rect 64 -181 84 -177
rect 788 -175 808 -171
rect 975 -175 995 -171
rect 788 -183 808 -179
rect 64 -189 84 -185
rect 975 -183 995 -179
rect 788 -191 808 -187
rect 975 -191 995 -187
rect 879 -197 899 -193
rect 879 -205 899 -201
rect 147 -232 151 -212
rect 155 -232 159 -212
rect 219 -217 239 -213
rect 219 -225 239 -221
rect 297 -225 301 -205
rect 305 -225 309 -205
rect 349 -225 369 -221
rect 64 -238 104 -234
rect 64 -246 104 -242
rect 219 -233 239 -229
rect 219 -241 239 -237
rect 349 -233 369 -229
rect 441 -234 445 -214
rect 449 -234 453 -214
rect 489 -219 509 -215
rect 489 -227 509 -223
rect 571 -225 575 -205
rect 579 -225 583 -205
rect 694 -225 698 -205
rect 702 -225 706 -205
rect 879 -213 899 -209
rect 349 -241 369 -237
rect 64 -254 104 -250
rect 219 -249 239 -245
rect 349 -249 369 -245
rect 219 -257 239 -253
rect 489 -235 509 -231
rect 489 -243 509 -239
rect 621 -230 641 -226
rect 621 -238 641 -234
rect 349 -257 369 -253
rect 621 -246 641 -242
rect 742 -246 842 -242
rect 742 -254 842 -250
rect 883 -253 887 -233
rect 891 -253 895 -233
rect 1040 -250 1060 -246
rect 742 -262 842 -258
rect 742 -270 842 -266
rect 1040 -258 1060 -254
rect 1040 -266 1060 -262
rect 742 -278 842 -274
rect 137 -300 141 -280
rect 145 -300 149 -280
rect 742 -286 842 -282
rect 949 -284 969 -280
rect 1136 -284 1156 -280
rect 949 -292 969 -288
rect 1136 -292 1156 -288
rect 949 -300 969 -296
rect 1136 -300 1156 -296
rect 64 -305 84 -301
rect 64 -313 84 -309
rect 1040 -306 1060 -302
rect 64 -321 84 -317
rect 257 -329 267 -325
rect 257 -337 267 -333
rect 147 -364 151 -344
rect 155 -364 159 -344
rect 257 -345 267 -341
rect 338 -344 342 -324
rect 346 -344 350 -324
rect 386 -325 406 -321
rect 386 -333 406 -329
rect 464 -333 468 -313
rect 472 -333 476 -313
rect 518 -324 538 -320
rect 518 -332 538 -328
rect 386 -341 406 -337
rect 257 -353 267 -349
rect 257 -361 267 -357
rect 64 -370 104 -366
rect 64 -378 104 -374
rect 386 -349 406 -345
rect 611 -333 615 -313
rect 619 -333 623 -313
rect 668 -327 688 -323
rect 518 -340 538 -336
rect 518 -348 538 -344
rect 386 -357 406 -353
rect 257 -369 267 -365
rect 668 -335 688 -331
rect 750 -333 754 -313
rect 758 -333 762 -313
rect 864 -333 868 -313
rect 872 -333 876 -313
rect 1040 -314 1060 -310
rect 1040 -322 1060 -318
rect 668 -343 688 -339
rect 518 -356 538 -352
rect 668 -351 688 -347
rect 791 -338 811 -334
rect 791 -346 811 -342
rect 791 -354 811 -350
rect 919 -359 1039 -355
rect 386 -365 406 -361
rect 919 -367 1039 -363
rect 257 -377 267 -373
rect 919 -375 1039 -371
rect 1089 -374 1093 -354
rect 1097 -374 1101 -354
rect 1247 -361 1267 -357
rect 1247 -369 1267 -365
rect 64 -386 104 -382
rect 919 -383 1039 -379
rect 919 -391 1039 -387
rect 1247 -377 1267 -373
rect 919 -399 1039 -395
rect 1156 -395 1176 -391
rect 1343 -395 1363 -391
rect 919 -407 1039 -403
rect 1156 -403 1176 -399
rect 1343 -403 1363 -399
rect 1156 -411 1176 -407
rect 1343 -411 1363 -407
rect 137 -433 141 -413
rect 145 -433 149 -413
rect 1247 -417 1267 -413
rect 1247 -425 1267 -421
rect 1247 -433 1267 -429
rect 64 -438 84 -434
rect 64 -446 84 -442
rect 64 -454 84 -450
rect 147 -497 151 -477
rect 155 -497 159 -477
rect 64 -503 104 -499
rect 64 -511 104 -507
rect 64 -519 104 -515
<< polysilicon >>
rect 142 116 144 119
rect 293 116 295 119
rect 55 88 64 90
rect 84 88 97 90
rect 117 88 120 90
rect 55 80 64 82
rect 84 80 97 82
rect 117 80 120 82
rect 142 80 144 96
rect 206 88 215 90
rect 235 88 248 90
rect 268 88 271 90
rect 206 80 215 82
rect 235 80 248 82
rect 268 80 271 82
rect 293 80 295 96
rect 460 76 472 78
rect 492 76 508 78
rect 528 76 531 78
rect 142 67 144 70
rect 293 67 295 70
rect 460 68 472 70
rect 492 68 508 70
rect 528 68 531 70
rect 152 52 154 55
rect 314 52 316 55
rect 369 42 381 44
rect 401 42 417 44
rect 437 42 440 44
rect 556 42 568 44
rect 588 42 604 44
rect 624 42 627 44
rect 369 34 381 36
rect 401 34 417 36
rect 437 34 440 36
rect 55 23 64 25
rect 104 23 116 25
rect 126 23 129 25
rect 55 15 64 17
rect 104 15 116 17
rect 126 15 129 17
rect 152 16 154 32
rect 217 23 226 25
rect 266 23 278 25
rect 288 23 291 25
rect 217 15 226 17
rect 266 15 278 17
rect 288 15 292 17
rect 314 16 316 32
rect 556 34 568 36
rect 588 34 604 36
rect 624 34 627 36
rect 460 20 472 22
rect 492 20 508 22
rect 528 20 531 22
rect 460 12 472 14
rect 492 12 508 14
rect 528 12 531 14
rect 152 3 154 6
rect 314 3 316 6
rect 142 -16 144 -13
rect 293 -16 295 -13
rect 414 -16 416 -13
rect 570 -16 572 -13
rect 197 -33 206 -31
rect 226 -33 238 -31
rect 268 -33 271 -31
rect 55 -44 64 -42
rect 84 -44 97 -42
rect 117 -44 120 -42
rect 55 -52 64 -50
rect 84 -52 97 -50
rect 117 -52 120 -50
rect 142 -52 144 -36
rect 454 -34 463 -32
rect 523 -34 535 -32
rect 545 -34 548 -32
rect 197 -41 206 -39
rect 226 -41 238 -39
rect 268 -41 271 -39
rect 197 -49 206 -47
rect 226 -49 238 -47
rect 268 -49 271 -47
rect 293 -52 295 -36
rect 327 -44 336 -42
rect 356 -44 369 -42
rect 389 -44 392 -42
rect 327 -52 336 -50
rect 356 -52 369 -50
rect 389 -52 392 -50
rect 414 -52 416 -36
rect 714 -34 726 -32
rect 746 -34 762 -32
rect 782 -34 785 -32
rect 454 -42 463 -40
rect 523 -42 535 -40
rect 545 -42 548 -40
rect 454 -50 463 -48
rect 523 -50 535 -48
rect 545 -50 548 -48
rect 570 -52 572 -36
rect 714 -42 726 -40
rect 746 -42 762 -40
rect 782 -42 785 -40
rect 142 -65 144 -62
rect 293 -65 295 -62
rect 414 -65 416 -62
rect 570 -65 572 -62
rect 623 -68 635 -66
rect 655 -68 671 -66
rect 691 -68 694 -66
rect 810 -68 822 -66
rect 842 -68 858 -66
rect 878 -68 881 -66
rect 623 -76 635 -74
rect 655 -76 671 -74
rect 691 -76 694 -74
rect 152 -80 154 -77
rect 810 -76 822 -74
rect 842 -76 858 -74
rect 878 -76 881 -74
rect 714 -90 726 -88
rect 746 -90 762 -88
rect 782 -90 785 -88
rect 313 -98 315 -95
rect 443 -98 445 -95
rect 560 -98 562 -95
rect 55 -109 64 -107
rect 104 -109 116 -107
rect 126 -109 129 -107
rect 55 -117 64 -115
rect 104 -117 116 -115
rect 126 -117 129 -115
rect 152 -116 154 -100
rect 207 -112 216 -110
rect 236 -112 248 -110
rect 288 -112 291 -110
rect 347 -115 356 -113
rect 376 -115 388 -113
rect 418 -115 421 -113
rect 207 -120 216 -118
rect 236 -120 248 -118
rect 288 -120 291 -118
rect 152 -129 154 -126
rect 207 -128 216 -126
rect 236 -128 248 -126
rect 288 -128 298 -126
rect 207 -136 216 -134
rect 236 -136 248 -134
rect 288 -136 291 -134
rect 296 -138 298 -128
rect 313 -134 315 -118
rect 714 -98 726 -96
rect 746 -98 762 -96
rect 782 -98 785 -96
rect 347 -123 356 -121
rect 376 -123 388 -121
rect 418 -123 421 -121
rect 347 -131 356 -129
rect 376 -131 388 -129
rect 418 -131 421 -129
rect 443 -134 445 -118
rect 473 -126 482 -124
rect 502 -126 515 -124
rect 535 -126 538 -124
rect 473 -134 482 -132
rect 502 -134 515 -132
rect 535 -134 538 -132
rect 560 -134 562 -118
rect 731 -127 733 -124
rect 594 -139 603 -137
rect 683 -139 695 -137
rect 705 -139 708 -137
rect 142 -148 144 -145
rect 313 -147 315 -144
rect 443 -147 445 -144
rect 560 -147 562 -144
rect 594 -147 603 -145
rect 683 -147 695 -145
rect 705 -147 708 -145
rect 867 -144 879 -142
rect 899 -144 915 -142
rect 935 -144 938 -142
rect 594 -155 603 -153
rect 683 -155 695 -153
rect 705 -155 708 -153
rect 594 -163 603 -161
rect 683 -163 695 -161
rect 705 -163 708 -161
rect 731 -163 733 -147
rect 867 -152 879 -150
rect 899 -152 915 -150
rect 935 -152 938 -150
rect 55 -176 64 -174
rect 84 -176 97 -174
rect 117 -176 120 -174
rect 55 -184 64 -182
rect 84 -184 97 -182
rect 117 -184 120 -182
rect 142 -184 144 -168
rect 731 -176 733 -173
rect 776 -178 788 -176
rect 808 -178 824 -176
rect 844 -178 847 -176
rect 963 -178 975 -176
rect 995 -178 1011 -176
rect 1031 -178 1034 -176
rect 776 -186 788 -184
rect 808 -186 824 -184
rect 844 -186 847 -184
rect 963 -186 975 -184
rect 995 -186 1011 -184
rect 1031 -186 1034 -184
rect 142 -197 144 -194
rect 867 -200 879 -198
rect 899 -200 915 -198
rect 935 -200 938 -198
rect 302 -205 304 -202
rect 576 -205 578 -202
rect 699 -205 701 -202
rect 152 -212 154 -209
rect 210 -220 219 -218
rect 239 -220 251 -218
rect 276 -220 279 -218
rect 446 -214 448 -211
rect 210 -228 219 -226
rect 239 -228 251 -226
rect 276 -228 279 -226
rect 55 -241 64 -239
rect 104 -241 116 -239
rect 126 -241 129 -239
rect 55 -249 64 -247
rect 104 -249 116 -247
rect 126 -249 129 -247
rect 152 -248 154 -232
rect 210 -236 219 -234
rect 239 -236 251 -234
rect 276 -236 282 -234
rect 302 -241 304 -225
rect 340 -228 349 -226
rect 369 -228 381 -226
rect 421 -228 424 -226
rect 480 -222 489 -220
rect 509 -222 521 -220
rect 551 -222 554 -220
rect 867 -208 879 -206
rect 899 -208 915 -206
rect 935 -208 938 -206
rect 480 -230 489 -228
rect 509 -230 521 -228
rect 551 -230 554 -228
rect 340 -236 349 -234
rect 369 -236 381 -234
rect 421 -236 424 -234
rect 210 -244 219 -242
rect 239 -244 251 -242
rect 276 -244 289 -242
rect 287 -248 289 -244
rect 210 -252 219 -250
rect 239 -252 251 -250
rect 276 -252 279 -250
rect 340 -244 349 -242
rect 369 -244 381 -242
rect 421 -244 424 -242
rect 302 -254 304 -251
rect 446 -250 448 -234
rect 480 -238 489 -236
rect 509 -238 521 -236
rect 551 -238 554 -236
rect 576 -241 578 -225
rect 612 -233 621 -231
rect 641 -233 654 -231
rect 674 -233 677 -231
rect 340 -252 349 -250
rect 369 -252 381 -250
rect 421 -252 424 -250
rect 152 -261 154 -258
rect 612 -241 621 -239
rect 641 -241 654 -239
rect 674 -241 677 -239
rect 699 -241 701 -225
rect 888 -233 890 -230
rect 733 -249 742 -247
rect 842 -249 854 -247
rect 864 -249 867 -247
rect 576 -254 578 -251
rect 699 -254 701 -251
rect 733 -257 742 -255
rect 842 -257 854 -255
rect 864 -257 867 -255
rect 446 -263 448 -260
rect 733 -265 742 -263
rect 842 -265 854 -263
rect 864 -265 867 -263
rect 888 -269 890 -253
rect 1028 -253 1040 -251
rect 1060 -253 1076 -251
rect 1096 -253 1099 -251
rect 1028 -261 1040 -259
rect 1060 -261 1076 -259
rect 1096 -261 1099 -259
rect 733 -273 742 -271
rect 842 -273 854 -271
rect 864 -273 867 -271
rect 142 -280 144 -277
rect 733 -281 742 -279
rect 842 -281 854 -279
rect 864 -281 867 -279
rect 888 -282 890 -279
rect 937 -287 949 -285
rect 969 -287 985 -285
rect 1005 -287 1008 -285
rect 1124 -287 1136 -285
rect 1156 -287 1172 -285
rect 1192 -287 1195 -285
rect 937 -295 949 -293
rect 969 -295 985 -293
rect 1005 -295 1008 -293
rect 1124 -295 1136 -293
rect 1156 -295 1172 -293
rect 1192 -295 1195 -293
rect 55 -308 64 -306
rect 84 -308 97 -306
rect 117 -308 120 -306
rect 55 -316 64 -314
rect 84 -316 97 -314
rect 117 -316 120 -314
rect 142 -316 144 -300
rect 1028 -309 1040 -307
rect 1060 -309 1076 -307
rect 1096 -309 1099 -307
rect 469 -313 471 -310
rect 616 -313 618 -310
rect 755 -313 757 -310
rect 869 -313 871 -310
rect 343 -324 345 -321
rect 142 -329 144 -326
rect 247 -332 257 -330
rect 267 -332 281 -330
rect 311 -332 314 -330
rect 247 -340 257 -338
rect 267 -340 281 -338
rect 311 -340 314 -338
rect 152 -344 154 -341
rect 377 -328 386 -326
rect 406 -328 418 -326
rect 443 -328 446 -326
rect 509 -327 518 -325
rect 538 -327 550 -325
rect 590 -327 593 -325
rect 377 -336 386 -334
rect 406 -336 418 -334
rect 443 -336 446 -334
rect 247 -348 257 -346
rect 267 -348 281 -346
rect 311 -348 314 -346
rect 247 -356 257 -354
rect 267 -356 281 -354
rect 311 -356 314 -354
rect 55 -373 64 -371
rect 104 -373 116 -371
rect 126 -373 129 -371
rect 55 -381 64 -379
rect 104 -381 116 -379
rect 126 -381 129 -379
rect 152 -380 154 -364
rect 343 -360 345 -344
rect 377 -344 386 -342
rect 406 -344 418 -342
rect 443 -344 446 -342
rect 469 -349 471 -333
rect 659 -330 668 -328
rect 688 -330 700 -328
rect 730 -330 733 -328
rect 509 -335 518 -333
rect 538 -335 550 -333
rect 590 -335 593 -333
rect 509 -343 518 -341
rect 538 -343 550 -341
rect 590 -343 593 -341
rect 377 -352 386 -350
rect 406 -352 418 -350
rect 443 -352 446 -350
rect 247 -364 257 -362
rect 267 -364 281 -362
rect 311 -364 314 -362
rect 377 -360 386 -358
rect 406 -360 418 -358
rect 443 -360 446 -358
rect 616 -349 618 -333
rect 1028 -317 1040 -315
rect 1060 -317 1076 -315
rect 1096 -317 1099 -315
rect 659 -338 668 -336
rect 688 -338 700 -336
rect 730 -338 733 -336
rect 659 -346 668 -344
rect 688 -346 700 -344
rect 730 -346 733 -344
rect 509 -351 518 -349
rect 538 -351 550 -349
rect 590 -351 593 -349
rect 755 -349 757 -333
rect 782 -341 791 -339
rect 811 -341 824 -339
rect 844 -341 847 -339
rect 782 -349 791 -347
rect 811 -349 824 -347
rect 844 -349 847 -347
rect 869 -349 871 -333
rect 1094 -354 1096 -351
rect 469 -362 471 -359
rect 616 -362 618 -359
rect 755 -362 757 -359
rect 869 -362 871 -359
rect 908 -362 919 -360
rect 1039 -362 1051 -360
rect 1061 -362 1064 -360
rect 247 -372 257 -370
rect 267 -372 281 -370
rect 311 -372 314 -370
rect 343 -373 345 -370
rect 908 -370 919 -368
rect 1039 -370 1051 -368
rect 1061 -370 1064 -368
rect 1235 -364 1247 -362
rect 1267 -364 1283 -362
rect 1303 -364 1306 -362
rect 1235 -372 1247 -370
rect 1267 -372 1283 -370
rect 1303 -372 1306 -370
rect 908 -378 919 -376
rect 1039 -378 1051 -376
rect 1061 -378 1064 -376
rect 908 -386 919 -384
rect 1039 -386 1051 -384
rect 1061 -386 1064 -384
rect 152 -393 154 -390
rect 1094 -390 1096 -374
rect 908 -394 919 -392
rect 1039 -394 1051 -392
rect 1061 -394 1064 -392
rect 1144 -398 1156 -396
rect 1176 -398 1192 -396
rect 1212 -398 1215 -396
rect 908 -402 919 -400
rect 1039 -402 1051 -400
rect 1061 -402 1064 -400
rect 1094 -403 1096 -400
rect 1331 -398 1343 -396
rect 1363 -398 1379 -396
rect 1399 -398 1402 -396
rect 1144 -406 1156 -404
rect 1176 -406 1192 -404
rect 1212 -406 1215 -404
rect 142 -413 144 -410
rect 1331 -406 1343 -404
rect 1363 -406 1379 -404
rect 1399 -406 1402 -404
rect 1235 -420 1247 -418
rect 1267 -420 1283 -418
rect 1303 -420 1306 -418
rect 1235 -428 1247 -426
rect 1267 -428 1283 -426
rect 1303 -428 1306 -426
rect 55 -441 64 -439
rect 84 -441 97 -439
rect 117 -441 120 -439
rect 55 -449 64 -447
rect 84 -449 97 -447
rect 117 -449 120 -447
rect 142 -449 144 -433
rect 142 -462 144 -459
rect 152 -477 154 -474
rect 55 -506 64 -504
rect 104 -506 116 -504
rect 126 -506 129 -504
rect 55 -514 64 -512
rect 104 -514 116 -512
rect 126 -514 129 -512
rect 152 -513 154 -497
rect 152 -526 154 -523
<< polycontact >>
rect 51 87 55 91
rect 51 79 55 83
rect 138 83 142 87
rect 202 87 206 91
rect 202 79 206 83
rect 289 83 293 87
rect 456 75 460 79
rect 456 67 460 71
rect 365 41 369 45
rect 365 33 369 37
rect 552 41 556 45
rect 51 22 55 26
rect 51 14 55 18
rect 148 19 152 23
rect 213 22 217 26
rect 213 14 217 18
rect 310 19 314 23
rect 552 33 556 37
rect 456 19 460 23
rect 456 11 460 15
rect 193 -34 197 -30
rect 51 -45 55 -41
rect 51 -53 55 -49
rect 138 -49 142 -45
rect 193 -42 197 -38
rect 450 -35 454 -31
rect 193 -50 197 -46
rect 289 -49 293 -45
rect 323 -45 327 -41
rect 323 -53 327 -49
rect 410 -49 414 -45
rect 450 -43 454 -39
rect 710 -35 714 -31
rect 450 -51 454 -47
rect 566 -49 570 -45
rect 710 -43 714 -39
rect 619 -69 623 -65
rect 619 -77 623 -73
rect 806 -69 810 -65
rect 806 -77 810 -73
rect 710 -91 714 -87
rect 51 -110 55 -106
rect 51 -118 55 -114
rect 148 -113 152 -109
rect 203 -113 207 -109
rect 203 -121 207 -117
rect 343 -116 347 -112
rect 203 -129 207 -125
rect 203 -137 207 -133
rect 309 -131 313 -127
rect 343 -124 347 -120
rect 421 -116 425 -112
rect 710 -99 714 -95
rect 343 -132 347 -128
rect 439 -131 443 -127
rect 469 -127 473 -123
rect 469 -135 473 -131
rect 538 -127 542 -123
rect 556 -131 560 -127
rect 590 -140 594 -136
rect 590 -148 594 -144
rect 863 -145 867 -141
rect 590 -156 594 -152
rect 590 -164 594 -160
rect 727 -160 731 -156
rect 863 -153 867 -149
rect 51 -177 55 -173
rect 51 -185 55 -181
rect 138 -181 142 -177
rect 772 -179 776 -175
rect 772 -187 776 -183
rect 959 -179 963 -175
rect 959 -187 963 -183
rect 863 -201 867 -197
rect 206 -221 210 -217
rect 206 -229 210 -225
rect 51 -242 55 -238
rect 51 -250 55 -246
rect 148 -245 152 -241
rect 206 -237 210 -233
rect 206 -245 210 -241
rect 282 -237 286 -233
rect 298 -238 302 -234
rect 336 -229 340 -225
rect 336 -237 340 -233
rect 476 -223 480 -219
rect 476 -231 480 -227
rect 554 -223 558 -219
rect 863 -209 867 -205
rect 206 -253 210 -249
rect 287 -252 291 -248
rect 336 -245 340 -241
rect 336 -253 340 -249
rect 424 -245 428 -241
rect 442 -247 446 -243
rect 476 -239 480 -235
rect 572 -238 576 -234
rect 608 -234 612 -230
rect 608 -242 612 -238
rect 677 -234 681 -230
rect 695 -238 699 -234
rect 677 -242 681 -238
rect 729 -250 733 -246
rect 729 -258 733 -254
rect 729 -266 733 -262
rect 729 -274 733 -270
rect 884 -266 888 -262
rect 1024 -254 1028 -250
rect 1024 -262 1028 -258
rect 729 -282 733 -278
rect 933 -288 937 -284
rect 933 -296 937 -292
rect 1120 -288 1124 -284
rect 1120 -296 1124 -292
rect 51 -309 55 -305
rect 51 -317 55 -313
rect 138 -313 142 -309
rect 1024 -310 1028 -306
rect 243 -333 247 -329
rect 243 -341 247 -337
rect 243 -349 247 -345
rect 373 -329 377 -325
rect 373 -337 377 -333
rect 505 -328 509 -324
rect 243 -357 247 -353
rect 314 -349 318 -345
rect 51 -374 55 -370
rect 51 -382 55 -378
rect 148 -377 152 -373
rect 243 -365 247 -361
rect 314 -357 318 -353
rect 339 -357 343 -353
rect 373 -345 377 -341
rect 373 -353 377 -349
rect 446 -345 450 -341
rect 465 -346 469 -342
rect 505 -336 509 -332
rect 655 -331 659 -327
rect 505 -344 509 -340
rect 243 -373 247 -369
rect 314 -366 318 -362
rect 373 -361 377 -357
rect 446 -353 450 -349
rect 505 -352 509 -348
rect 593 -344 597 -340
rect 612 -346 616 -342
rect 655 -339 659 -335
rect 1024 -318 1028 -314
rect 655 -347 659 -343
rect 751 -346 755 -342
rect 593 -353 597 -349
rect 778 -342 782 -338
rect 778 -350 782 -346
rect 865 -346 869 -342
rect 904 -363 908 -359
rect 904 -371 908 -367
rect 904 -379 908 -375
rect 1231 -365 1235 -361
rect 1231 -373 1235 -369
rect 904 -387 908 -383
rect 904 -395 908 -391
rect 1090 -387 1094 -383
rect 904 -403 908 -399
rect 1140 -399 1144 -395
rect 1140 -407 1144 -403
rect 1327 -399 1331 -395
rect 1327 -407 1331 -403
rect 1231 -421 1235 -417
rect 1231 -429 1235 -425
rect 51 -442 55 -438
rect 51 -450 55 -446
rect 138 -446 142 -442
rect 51 -507 55 -503
rect 51 -515 55 -511
rect 148 -510 152 -506
<< metal1 >>
rect -1 138 8 144
rect -1 135 185 138
rect -1 119 173 122
rect 0 91 9 97
rect 0 88 30 91
rect 0 74 9 83
rect 19 16 22 88
rect 25 27 28 78
rect 19 13 25 16
rect 33 0 36 63
rect 39 58 42 119
rect 58 95 61 119
rect 137 116 141 119
rect 90 98 130 102
rect 90 95 94 98
rect 58 91 64 95
rect 90 91 97 95
rect 50 87 51 91
rect 50 79 51 83
rect 58 79 61 91
rect 90 87 94 91
rect 126 87 130 98
rect 145 87 149 96
rect 182 91 185 135
rect 198 119 352 122
rect 209 95 212 119
rect 288 116 292 119
rect 241 98 281 102
rect 241 95 245 98
rect 209 91 215 95
rect 241 91 248 95
rect 182 87 202 91
rect 84 83 94 87
rect 126 83 138 87
rect 145 83 175 87
rect 145 80 149 83
rect 58 75 64 79
rect 117 75 123 79
rect 120 67 123 75
rect 137 67 141 70
rect 51 64 141 67
rect 39 55 162 58
rect 39 9 42 55
rect 50 22 51 26
rect 50 14 51 18
rect 58 14 61 55
rect 147 52 151 55
rect 110 33 138 36
rect 110 30 113 33
rect 104 26 113 30
rect 110 22 113 26
rect 135 23 138 33
rect 171 46 175 83
rect 182 79 202 83
rect 209 79 212 91
rect 241 87 245 91
rect 277 87 281 98
rect 349 101 352 119
rect 349 97 562 101
rect 296 87 300 96
rect 235 83 245 87
rect 277 83 289 87
rect 296 83 313 87
rect 500 86 543 90
rect 296 80 300 83
rect 155 23 159 32
rect 182 23 186 79
rect 209 75 215 79
rect 268 75 274 79
rect 271 67 274 75
rect 288 67 292 70
rect 110 18 116 22
rect 135 19 148 23
rect 155 19 186 23
rect 191 64 292 67
rect 309 69 313 83
rect 463 79 472 83
rect 361 75 456 79
rect 155 16 159 19
rect 58 10 64 14
rect 126 10 132 14
rect 129 0 132 10
rect 147 0 151 6
rect 191 3 194 64
rect 202 55 313 58
rect 202 41 207 45
rect 203 18 207 41
rect 213 26 217 45
rect 203 14 213 18
rect 220 14 223 55
rect 309 52 313 55
rect 272 33 300 36
rect 272 30 275 33
rect 266 26 275 30
rect 288 26 294 30
rect 272 22 275 26
rect 272 18 278 22
rect 291 14 294 26
rect 297 23 300 33
rect 361 45 365 75
rect 452 56 456 71
rect 463 67 466 79
rect 500 75 504 86
rect 528 79 531 83
rect 492 71 504 75
rect 500 67 504 71
rect 409 52 456 56
rect 372 45 381 49
rect 332 41 365 45
rect 332 36 336 41
rect 317 23 321 32
rect 343 33 365 37
rect 372 33 375 45
rect 409 41 413 52
rect 437 45 441 49
rect 401 37 413 41
rect 409 33 413 37
rect 343 23 347 33
rect 297 19 310 23
rect 317 19 347 23
rect 317 16 321 19
rect 220 10 226 14
rect 288 10 294 14
rect 291 3 294 10
rect 361 15 365 33
rect 372 29 381 33
rect 409 29 417 33
rect 452 19 456 52
rect 463 63 472 67
rect 500 63 508 67
rect 463 54 467 63
rect 463 50 512 54
rect 463 27 467 50
rect 539 45 543 86
rect 558 54 562 97
rect 596 53 646 57
rect 559 45 568 49
rect 539 41 552 45
rect 539 34 552 37
rect 500 33 552 34
rect 559 33 562 45
rect 596 41 600 53
rect 624 45 628 49
rect 588 37 600 41
rect 596 33 600 37
rect 500 30 543 33
rect 463 23 472 27
rect 361 11 456 15
rect 463 11 466 23
rect 500 19 504 30
rect 559 29 568 33
rect 596 29 604 33
rect 528 23 538 27
rect 492 15 504 19
rect 500 11 504 15
rect 463 7 472 11
rect 500 7 508 11
rect 309 3 313 6
rect 534 4 538 23
rect 628 4 632 45
rect 349 3 632 4
rect 191 0 632 3
rect 33 -2 194 0
rect 33 -3 127 -2
rect 39 -11 41 -10
rect 132 -3 194 -2
rect 555 -10 816 -9
rect 46 -11 816 -10
rect 39 -13 816 -11
rect 0 -41 9 -35
rect 0 -44 30 -41
rect 0 -58 9 -49
rect 19 -116 22 -44
rect 25 -105 28 -54
rect 19 -119 25 -116
rect 33 -131 36 -69
rect 39 -74 42 -13
rect 58 -37 61 -13
rect 137 -16 141 -13
rect 90 -34 130 -30
rect 90 -37 94 -34
rect 58 -41 64 -37
rect 90 -41 97 -37
rect 50 -45 51 -41
rect 50 -53 51 -49
rect 58 -53 61 -41
rect 90 -45 94 -41
rect 126 -45 130 -34
rect 145 -45 149 -36
rect 178 -38 182 -21
rect 191 -30 193 -29
rect 188 -34 193 -30
rect 200 -34 203 -13
rect 288 -16 292 -13
rect 232 -23 282 -20
rect 232 -26 235 -23
rect 226 -30 238 -26
rect 200 -38 206 -34
rect 178 -42 193 -38
rect 84 -49 94 -45
rect 126 -49 138 -45
rect 145 -49 165 -45
rect 145 -52 149 -49
rect 173 -50 193 -46
rect 200 -50 203 -38
rect 231 -42 235 -30
rect 226 -46 235 -42
rect 271 -50 274 -26
rect 279 -45 282 -23
rect 296 -45 300 -36
rect 319 -45 323 -22
rect 330 -37 333 -13
rect 409 -16 413 -13
rect 362 -34 403 -30
rect 362 -37 366 -34
rect 330 -41 336 -37
rect 362 -41 369 -37
rect 279 -49 289 -45
rect 296 -49 306 -45
rect 58 -57 64 -53
rect 117 -57 123 -53
rect 120 -65 123 -57
rect 173 -57 177 -50
rect 200 -54 206 -50
rect 268 -54 274 -50
rect 296 -52 300 -49
rect 137 -65 141 -62
rect 271 -65 274 -54
rect 319 -57 323 -49
rect 330 -53 333 -41
rect 362 -45 366 -41
rect 400 -45 403 -34
rect 417 -45 421 -36
rect 432 -35 450 -31
rect 432 -45 436 -35
rect 356 -49 366 -45
rect 400 -49 410 -45
rect 417 -49 436 -45
rect 439 -43 450 -39
rect 417 -52 421 -49
rect 330 -57 336 -53
rect 389 -57 395 -53
rect 288 -65 292 -62
rect 392 -65 395 -57
rect 439 -57 443 -43
rect 447 -51 450 -47
rect 457 -51 460 -13
rect 565 -16 569 -13
rect 529 -24 559 -21
rect 529 -27 532 -24
rect 523 -31 535 -27
rect 529 -43 532 -31
rect 548 -35 551 -27
rect 545 -39 551 -35
rect 529 -47 535 -43
rect 548 -51 551 -39
rect 556 -45 559 -24
rect 573 -45 577 -36
rect 556 -49 566 -45
rect 573 -49 583 -45
rect 457 -55 463 -51
rect 545 -55 551 -51
rect 573 -52 577 -49
rect 457 -61 460 -55
rect 409 -65 413 -62
rect 548 -65 551 -55
rect 565 -65 569 -62
rect 51 -68 569 -65
rect 39 -77 151 -74
rect 311 -75 439 -72
rect 39 -123 42 -77
rect 50 -110 51 -106
rect 50 -118 51 -114
rect 58 -118 61 -77
rect 147 -80 151 -77
rect 110 -99 138 -96
rect 110 -102 113 -99
rect 104 -106 113 -102
rect 110 -110 113 -106
rect 135 -109 138 -99
rect 155 -109 159 -100
rect 184 -80 187 -76
rect 449 -80 452 -76
rect 184 -83 452 -80
rect 173 -109 177 -84
rect 185 -95 559 -92
rect 196 -109 201 -108
rect 210 -105 213 -95
rect 308 -98 312 -95
rect 242 -102 302 -99
rect 242 -105 245 -102
rect 210 -109 216 -105
rect 241 -109 248 -105
rect 110 -114 116 -110
rect 135 -113 148 -109
rect 155 -113 186 -109
rect 196 -113 203 -109
rect 155 -116 159 -113
rect 58 -122 64 -118
rect 126 -122 132 -118
rect 129 -131 132 -122
rect 182 -125 186 -113
rect 194 -121 203 -117
rect 210 -121 213 -109
rect 241 -113 245 -109
rect 236 -117 245 -113
rect 210 -125 216 -121
rect 147 -131 151 -126
rect 182 -129 203 -125
rect 33 -134 179 -131
rect 44 -144 141 -142
rect 39 -145 141 -144
rect 0 -173 9 -167
rect 0 -176 30 -173
rect 0 -190 9 -181
rect 19 -248 22 -176
rect 25 -237 28 -186
rect 19 -251 25 -248
rect 33 -264 36 -201
rect 39 -206 42 -145
rect 58 -169 61 -145
rect 137 -148 141 -145
rect 176 -147 179 -134
rect 184 -137 203 -133
rect 210 -137 213 -125
rect 241 -129 245 -117
rect 299 -127 302 -102
rect 339 -116 343 -112
rect 350 -116 353 -95
rect 438 -98 442 -95
rect 382 -105 432 -102
rect 382 -108 385 -105
rect 376 -112 388 -108
rect 316 -126 320 -118
rect 350 -120 356 -116
rect 339 -124 343 -120
rect 236 -133 245 -129
rect 299 -131 309 -127
rect 316 -134 320 -131
rect 184 -139 188 -137
rect 210 -141 216 -137
rect 288 -141 294 -137
rect 210 -144 213 -141
rect 291 -147 294 -141
rect 334 -132 343 -128
rect 350 -132 353 -120
rect 381 -124 385 -112
rect 376 -128 385 -124
rect 429 -127 432 -105
rect 446 -127 450 -118
rect 465 -127 469 -112
rect 476 -119 479 -95
rect 555 -98 559 -95
rect 565 -98 569 -68
rect 597 -65 601 -23
rect 754 -24 797 -20
rect 717 -31 726 -27
rect 615 -35 710 -31
rect 615 -65 619 -35
rect 706 -54 710 -39
rect 717 -43 720 -31
rect 754 -35 758 -24
rect 782 -31 785 -27
rect 746 -39 758 -35
rect 754 -43 758 -39
rect 663 -58 710 -54
rect 626 -65 635 -61
rect 597 -69 619 -65
rect 582 -77 619 -73
rect 626 -77 629 -65
rect 663 -69 667 -58
rect 691 -65 695 -61
rect 655 -73 667 -69
rect 663 -77 667 -73
rect 508 -116 552 -112
rect 508 -119 512 -116
rect 476 -123 482 -119
rect 508 -123 515 -119
rect 429 -131 439 -127
rect 446 -131 456 -127
rect 334 -139 338 -132
rect 350 -136 356 -132
rect 418 -136 424 -132
rect 446 -134 450 -131
rect 308 -147 312 -144
rect 421 -147 424 -136
rect 465 -139 469 -131
rect 476 -135 479 -123
rect 508 -127 512 -123
rect 548 -127 552 -116
rect 567 -106 569 -98
rect 615 -95 619 -77
rect 626 -81 635 -77
rect 663 -81 671 -77
rect 706 -91 710 -58
rect 717 -47 726 -43
rect 754 -47 762 -43
rect 717 -56 721 -47
rect 717 -60 766 -56
rect 717 -83 721 -60
rect 793 -65 797 -24
rect 812 -56 816 -13
rect 850 -57 900 -53
rect 813 -65 822 -61
rect 793 -69 806 -65
rect 793 -76 806 -73
rect 754 -77 806 -76
rect 813 -77 816 -65
rect 850 -69 854 -57
rect 878 -65 882 -61
rect 842 -73 854 -69
rect 850 -77 854 -73
rect 754 -80 797 -77
rect 717 -87 726 -83
rect 615 -99 710 -95
rect 717 -99 720 -87
rect 754 -91 758 -80
rect 813 -81 822 -77
rect 850 -81 858 -77
rect 782 -87 792 -83
rect 746 -95 758 -91
rect 754 -99 758 -95
rect 717 -103 726 -99
rect 754 -103 762 -99
rect 788 -106 792 -87
rect 882 -106 886 -65
rect 567 -110 886 -106
rect 563 -127 567 -118
rect 723 -120 969 -119
rect 585 -123 969 -120
rect 502 -131 512 -127
rect 548 -131 556 -127
rect 563 -131 579 -127
rect 563 -134 567 -131
rect 476 -139 482 -135
rect 535 -139 541 -135
rect 438 -147 442 -144
rect 538 -147 541 -139
rect 575 -136 579 -131
rect 575 -140 590 -136
rect 555 -147 559 -144
rect 90 -166 130 -162
rect 90 -169 94 -166
rect 58 -173 64 -169
rect 90 -173 97 -169
rect 50 -177 51 -173
rect 50 -185 51 -181
rect 58 -185 61 -173
rect 90 -177 94 -173
rect 126 -177 130 -166
rect 176 -150 559 -147
rect 461 -157 543 -154
rect 145 -177 149 -168
rect 84 -181 94 -177
rect 126 -181 138 -177
rect 145 -181 165 -177
rect 145 -184 149 -181
rect 58 -189 64 -185
rect 117 -189 123 -185
rect 120 -197 123 -189
rect 179 -186 183 -168
rect 302 -178 305 -160
rect 426 -164 429 -158
rect 327 -167 429 -164
rect 327 -178 330 -167
rect 480 -178 483 -166
rect 555 -176 559 -150
rect 570 -148 590 -144
rect 570 -158 574 -148
rect 577 -156 590 -152
rect 577 -162 581 -156
rect 573 -166 581 -162
rect 586 -168 590 -160
rect 597 -164 600 -123
rect 688 -129 720 -126
rect 688 -132 691 -129
rect 683 -136 691 -132
rect 705 -136 711 -132
rect 687 -140 691 -136
rect 687 -144 695 -140
rect 687 -156 691 -144
rect 708 -148 711 -136
rect 705 -152 711 -148
rect 687 -160 695 -156
rect 708 -164 711 -152
rect 717 -156 720 -129
rect 726 -127 730 -123
rect 907 -134 950 -130
rect 870 -141 879 -137
rect 734 -156 738 -147
rect 768 -145 863 -141
rect 717 -160 727 -156
rect 734 -160 742 -156
rect 734 -163 738 -160
rect 597 -168 603 -164
rect 705 -168 711 -164
rect 708 -176 711 -168
rect 726 -176 730 -173
rect 768 -175 772 -145
rect 859 -164 863 -149
rect 870 -153 873 -141
rect 907 -145 911 -134
rect 935 -141 938 -137
rect 899 -149 911 -145
rect 907 -153 911 -149
rect 816 -168 863 -164
rect 779 -175 788 -171
rect 555 -179 730 -176
rect 179 -187 706 -186
rect 165 -190 706 -187
rect 165 -191 183 -190
rect 137 -197 141 -194
rect 51 -200 141 -197
rect 147 -202 157 -198
rect 147 -206 151 -202
rect 39 -209 151 -206
rect 165 -205 169 -191
rect 177 -199 183 -197
rect 177 -200 721 -199
rect 180 -202 721 -200
rect 165 -209 183 -205
rect 39 -255 42 -209
rect 50 -242 51 -238
rect 50 -250 51 -246
rect 58 -250 61 -209
rect 147 -212 151 -209
rect 110 -231 138 -228
rect 110 -234 113 -231
rect 104 -238 113 -234
rect 110 -242 113 -238
rect 135 -241 138 -231
rect 155 -241 159 -232
rect 179 -241 183 -209
rect 197 -209 201 -205
rect 202 -221 206 -210
rect 213 -221 216 -202
rect 297 -205 301 -202
rect 245 -210 292 -207
rect 245 -213 248 -210
rect 239 -217 251 -213
rect 192 -225 196 -221
rect 213 -225 219 -221
rect 192 -229 206 -225
rect 193 -237 206 -233
rect 213 -237 216 -225
rect 244 -229 248 -217
rect 239 -233 248 -229
rect 213 -241 219 -237
rect 110 -246 116 -242
rect 135 -245 148 -241
rect 155 -245 206 -241
rect 155 -248 159 -245
rect 58 -254 64 -250
rect 126 -254 132 -250
rect 129 -264 132 -254
rect 172 -249 176 -245
rect 191 -253 206 -249
rect 213 -253 216 -241
rect 244 -245 248 -233
rect 289 -234 292 -210
rect 343 -208 346 -202
rect 343 -211 459 -208
rect 331 -217 336 -212
rect 305 -234 309 -225
rect 333 -229 336 -217
rect 343 -221 346 -211
rect 441 -214 445 -211
rect 375 -218 438 -215
rect 375 -221 378 -218
rect 343 -225 349 -221
rect 374 -225 381 -221
rect 326 -233 330 -229
rect 289 -238 298 -234
rect 305 -238 318 -234
rect 326 -237 336 -233
rect 343 -237 346 -225
rect 374 -229 378 -225
rect 369 -233 378 -229
rect 305 -241 309 -238
rect 239 -249 248 -245
rect 314 -246 318 -238
rect 343 -241 349 -237
rect 324 -244 336 -241
rect 329 -245 336 -244
rect 191 -254 196 -253
rect 147 -264 151 -258
rect 213 -257 219 -253
rect 276 -257 282 -253
rect 279 -263 282 -257
rect 297 -263 301 -251
rect 332 -253 336 -249
rect 343 -253 346 -241
rect 374 -245 378 -233
rect 435 -243 438 -218
rect 472 -223 476 -212
rect 483 -223 486 -202
rect 571 -205 575 -202
rect 515 -212 565 -209
rect 515 -215 518 -212
rect 509 -219 521 -215
rect 460 -227 464 -224
rect 483 -227 489 -223
rect 460 -231 476 -227
rect 449 -243 453 -234
rect 469 -239 476 -235
rect 483 -239 486 -227
rect 514 -231 518 -219
rect 509 -235 518 -231
rect 562 -234 565 -212
rect 605 -217 608 -212
rect 579 -234 583 -225
rect 604 -234 608 -217
rect 615 -226 618 -202
rect 694 -205 698 -202
rect 647 -222 688 -219
rect 647 -226 651 -222
rect 615 -230 621 -226
rect 647 -230 654 -226
rect 562 -238 572 -234
rect 579 -238 589 -234
rect 369 -249 378 -245
rect 435 -247 442 -243
rect 449 -247 463 -243
rect 449 -250 453 -247
rect 343 -257 349 -253
rect 421 -257 427 -253
rect 343 -260 346 -257
rect 424 -263 427 -257
rect 459 -253 463 -247
rect 469 -245 473 -239
rect 483 -243 489 -239
rect 551 -243 557 -239
rect 579 -241 583 -238
rect 554 -254 557 -243
rect 604 -246 608 -238
rect 615 -242 618 -230
rect 647 -234 651 -230
rect 685 -234 688 -222
rect 702 -234 706 -225
rect 718 -227 721 -202
rect 726 -216 730 -179
rect 741 -179 772 -175
rect 741 -186 745 -179
rect 738 -190 745 -186
rect 756 -187 772 -183
rect 779 -187 782 -175
rect 816 -179 820 -168
rect 844 -175 848 -171
rect 808 -183 820 -179
rect 816 -187 820 -183
rect 768 -205 772 -187
rect 779 -191 788 -187
rect 816 -191 824 -187
rect 859 -201 863 -168
rect 870 -157 879 -153
rect 907 -157 915 -153
rect 870 -166 874 -157
rect 870 -170 919 -166
rect 870 -193 874 -170
rect 946 -175 950 -134
rect 965 -166 969 -123
rect 1003 -167 1053 -163
rect 966 -175 975 -171
rect 946 -179 959 -175
rect 946 -186 959 -183
rect 907 -187 959 -186
rect 966 -187 969 -175
rect 1003 -179 1007 -167
rect 1031 -175 1035 -171
rect 995 -183 1007 -179
rect 1003 -187 1007 -183
rect 907 -190 950 -187
rect 870 -197 879 -193
rect 768 -209 863 -205
rect 870 -209 873 -197
rect 907 -201 911 -190
rect 966 -191 975 -187
rect 1003 -191 1011 -187
rect 935 -197 945 -193
rect 899 -205 911 -201
rect 907 -209 911 -205
rect 870 -213 879 -209
rect 907 -213 915 -209
rect 941 -216 945 -197
rect 1035 -216 1039 -175
rect 726 -220 1039 -216
rect 718 -228 921 -227
rect 718 -230 1130 -228
rect 641 -238 651 -234
rect 685 -238 695 -234
rect 702 -238 729 -234
rect 702 -241 706 -238
rect 615 -246 621 -242
rect 604 -251 605 -246
rect 571 -254 575 -251
rect 651 -254 654 -242
rect 725 -250 729 -238
rect 694 -254 698 -251
rect 472 -257 698 -254
rect 441 -263 445 -260
rect 472 -263 475 -257
rect 160 -264 475 -263
rect 33 -266 475 -264
rect 33 -267 127 -266
rect 132 -267 163 -266
rect 39 -276 40 -274
rect 45 -276 141 -274
rect 39 -277 141 -276
rect 0 -305 9 -299
rect 0 -308 30 -305
rect 0 -322 9 -313
rect 19 -380 22 -308
rect 25 -369 28 -318
rect 19 -383 25 -380
rect 33 -396 36 -333
rect 39 -338 42 -277
rect 58 -301 61 -277
rect 137 -280 141 -277
rect 90 -298 130 -294
rect 90 -301 94 -298
rect 58 -305 64 -301
rect 90 -305 97 -301
rect 50 -309 51 -305
rect 50 -317 51 -313
rect 58 -317 61 -305
rect 90 -309 94 -305
rect 126 -309 130 -298
rect 187 -281 192 -280
rect 187 -285 196 -281
rect 145 -309 149 -300
rect 84 -313 94 -309
rect 126 -313 138 -309
rect 145 -313 178 -309
rect 145 -316 149 -313
rect 58 -321 64 -317
rect 117 -321 123 -317
rect 120 -329 123 -321
rect 137 -329 141 -326
rect 51 -332 141 -329
rect 39 -341 165 -338
rect 39 -387 42 -341
rect 50 -374 51 -370
rect 50 -382 51 -378
rect 58 -382 61 -341
rect 147 -344 151 -341
rect 110 -363 138 -360
rect 110 -366 113 -363
rect 104 -370 113 -366
rect 110 -374 113 -370
rect 135 -373 138 -363
rect 155 -373 159 -364
rect 192 -364 196 -285
rect 204 -289 207 -274
rect 204 -292 242 -289
rect 206 -345 210 -325
rect 227 -337 231 -307
rect 239 -329 242 -292
rect 262 -301 265 -274
rect 280 -293 283 -274
rect 694 -296 698 -257
rect 707 -258 729 -254
rect 703 -266 729 -262
rect 703 -272 707 -266
rect 713 -274 729 -270
rect 713 -282 717 -274
rect 707 -286 717 -282
rect 722 -282 729 -278
rect 736 -282 739 -230
rect 883 -233 887 -230
rect 917 -232 1130 -230
rect 848 -239 877 -236
rect 848 -242 851 -239
rect 842 -246 854 -242
rect 847 -258 851 -246
rect 864 -254 870 -250
rect 847 -262 854 -258
rect 847 -274 851 -262
rect 867 -266 870 -254
rect 874 -262 877 -239
rect 1068 -243 1111 -239
rect 1031 -250 1040 -246
rect 891 -262 895 -253
rect 929 -254 1024 -250
rect 874 -266 884 -262
rect 891 -266 901 -262
rect 864 -270 870 -266
rect 891 -269 895 -266
rect 847 -278 854 -274
rect 867 -282 870 -270
rect 722 -286 726 -282
rect 736 -286 742 -282
rect 864 -283 870 -282
rect 883 -283 887 -279
rect 864 -286 887 -283
rect 917 -284 921 -271
rect 929 -284 933 -254
rect 1020 -273 1024 -258
rect 1031 -262 1034 -250
rect 1068 -254 1072 -243
rect 1096 -250 1099 -246
rect 1060 -258 1072 -254
rect 1068 -262 1072 -258
rect 977 -277 1024 -273
rect 940 -284 949 -280
rect 736 -292 739 -286
rect 867 -296 870 -286
rect 694 -299 870 -296
rect 262 -304 362 -301
rect 250 -310 868 -307
rect 250 -325 254 -310
rect 273 -322 335 -318
rect 273 -325 277 -322
rect 250 -329 257 -325
rect 273 -329 281 -325
rect 239 -333 243 -329
rect 227 -341 243 -337
rect 250 -341 254 -329
rect 273 -333 277 -329
rect 267 -337 277 -333
rect 250 -345 257 -341
rect 206 -349 243 -345
rect 208 -354 243 -353
rect 213 -357 243 -354
rect 250 -357 254 -345
rect 273 -349 277 -337
rect 267 -353 277 -349
rect 331 -353 335 -322
rect 338 -324 342 -310
rect 369 -329 373 -319
rect 380 -329 383 -310
rect 464 -313 468 -310
rect 412 -318 461 -315
rect 412 -321 415 -318
rect 406 -325 418 -321
rect 380 -333 386 -329
rect 360 -337 373 -333
rect 346 -353 350 -344
rect 360 -345 373 -341
rect 380 -345 383 -333
rect 411 -337 415 -325
rect 406 -341 415 -337
rect 360 -352 363 -345
rect 380 -349 386 -345
rect 250 -361 257 -357
rect 217 -364 243 -361
rect 192 -365 243 -364
rect 192 -368 221 -365
rect 192 -373 196 -368
rect 110 -378 116 -374
rect 135 -377 148 -373
rect 155 -377 196 -373
rect 239 -377 243 -369
rect 250 -373 254 -361
rect 273 -365 277 -353
rect 331 -357 339 -353
rect 346 -357 356 -353
rect 346 -360 350 -357
rect 267 -369 277 -365
rect 338 -373 342 -370
rect 155 -380 159 -377
rect 58 -386 64 -382
rect 126 -386 132 -382
rect 129 -396 132 -386
rect 201 -381 243 -377
rect 250 -377 257 -373
rect 311 -377 342 -373
rect 147 -396 151 -390
rect 33 -399 159 -396
rect 39 -409 40 -407
rect 45 -409 177 -407
rect 39 -410 177 -409
rect 0 -438 9 -432
rect 0 -441 30 -438
rect 0 -455 9 -446
rect 19 -513 22 -441
rect 25 -502 28 -451
rect 19 -516 25 -513
rect 33 -529 36 -466
rect 39 -471 42 -410
rect 58 -434 61 -410
rect 137 -413 141 -410
rect 90 -431 130 -427
rect 90 -434 94 -431
rect 58 -438 64 -434
rect 90 -438 97 -434
rect 50 -442 51 -438
rect 50 -450 51 -446
rect 58 -450 61 -438
rect 90 -442 94 -438
rect 126 -442 130 -431
rect 145 -442 149 -433
rect 201 -419 205 -381
rect 250 -407 254 -377
rect 338 -391 342 -377
rect 380 -361 383 -349
rect 411 -353 415 -341
rect 458 -342 461 -318
rect 503 -318 505 -313
rect 501 -328 505 -318
rect 512 -320 515 -310
rect 611 -313 615 -310
rect 544 -317 608 -314
rect 544 -320 547 -317
rect 512 -324 518 -320
rect 543 -324 550 -320
rect 458 -346 465 -342
rect 472 -349 476 -333
rect 490 -335 505 -332
rect 485 -336 505 -335
rect 512 -336 515 -324
rect 543 -328 547 -324
rect 538 -332 547 -328
rect 512 -340 518 -336
rect 483 -342 505 -340
rect 488 -344 505 -342
rect 406 -357 415 -353
rect 501 -352 505 -348
rect 512 -352 515 -340
rect 543 -344 547 -332
rect 605 -342 608 -317
rect 647 -321 655 -317
rect 651 -331 655 -321
rect 662 -331 665 -310
rect 750 -313 754 -310
rect 694 -320 744 -317
rect 694 -323 697 -320
rect 688 -327 700 -323
rect 619 -342 623 -333
rect 638 -335 641 -334
rect 662 -335 668 -331
rect 638 -339 655 -335
rect 538 -348 547 -344
rect 605 -346 612 -342
rect 619 -346 629 -342
rect 512 -356 518 -352
rect 548 -356 550 -352
rect 619 -349 623 -346
rect 651 -348 655 -343
rect 662 -347 665 -335
rect 693 -339 697 -327
rect 688 -343 697 -339
rect 741 -342 744 -320
rect 758 -342 762 -333
rect 785 -334 788 -310
rect 864 -313 868 -310
rect 817 -331 857 -327
rect 817 -334 821 -331
rect 785 -338 791 -334
rect 817 -338 824 -334
rect 773 -342 778 -338
rect 741 -346 751 -342
rect 758 -346 765 -342
rect 512 -359 515 -356
rect 380 -365 386 -361
rect 443 -362 446 -361
rect 443 -365 449 -362
rect 346 -376 350 -370
rect 446 -371 449 -365
rect 464 -370 468 -359
rect 548 -362 551 -356
rect 654 -353 655 -348
rect 662 -351 668 -347
rect 730 -351 736 -347
rect 758 -349 762 -346
rect 611 -362 615 -359
rect 733 -362 736 -351
rect 774 -350 778 -346
rect 785 -350 788 -338
rect 817 -342 821 -338
rect 853 -342 857 -331
rect 883 -325 887 -286
rect 917 -288 933 -284
rect 906 -292 911 -290
rect 906 -296 933 -292
rect 940 -296 943 -284
rect 977 -288 981 -277
rect 1005 -284 1009 -280
rect 969 -292 981 -288
rect 977 -296 981 -292
rect 929 -314 933 -296
rect 940 -300 949 -296
rect 977 -300 985 -296
rect 1020 -310 1024 -277
rect 1031 -266 1040 -262
rect 1068 -266 1076 -262
rect 1031 -275 1035 -266
rect 1031 -279 1080 -275
rect 1031 -302 1035 -279
rect 1107 -284 1111 -243
rect 1126 -275 1130 -232
rect 1164 -276 1214 -272
rect 1127 -284 1136 -280
rect 1107 -288 1120 -284
rect 1107 -295 1120 -292
rect 1068 -296 1120 -295
rect 1127 -296 1130 -284
rect 1164 -288 1168 -276
rect 1192 -284 1196 -280
rect 1156 -292 1168 -288
rect 1164 -296 1168 -292
rect 1068 -299 1111 -296
rect 1031 -306 1040 -302
rect 929 -318 1024 -314
rect 1031 -318 1034 -306
rect 1068 -310 1072 -299
rect 1127 -300 1136 -296
rect 1164 -300 1172 -296
rect 1096 -306 1106 -302
rect 1060 -314 1072 -310
rect 1068 -318 1072 -314
rect 1031 -322 1040 -318
rect 1068 -322 1076 -318
rect 1102 -325 1106 -306
rect 1196 -325 1200 -284
rect 883 -329 1200 -325
rect 872 -342 876 -333
rect 811 -346 821 -342
rect 853 -346 865 -342
rect 872 -346 904 -342
rect 872 -349 876 -346
rect 785 -354 791 -350
rect 844 -354 850 -350
rect 750 -362 754 -359
rect 847 -362 850 -354
rect 864 -362 868 -359
rect 501 -365 868 -362
rect 900 -363 904 -346
rect 911 -343 1337 -339
rect 501 -370 504 -365
rect 464 -371 504 -370
rect 369 -374 504 -371
rect 346 -380 358 -376
rect 369 -391 372 -374
rect 215 -411 254 -407
rect 259 -395 372 -391
rect 201 -423 245 -419
rect 84 -446 94 -442
rect 126 -446 138 -442
rect 145 -446 180 -442
rect 145 -449 149 -446
rect 58 -454 64 -450
rect 117 -454 123 -450
rect 120 -462 123 -454
rect 137 -462 141 -459
rect 51 -465 141 -462
rect 39 -474 165 -471
rect 39 -520 42 -474
rect 50 -507 51 -503
rect 50 -515 51 -511
rect 58 -515 61 -474
rect 147 -477 151 -474
rect 110 -496 138 -493
rect 110 -499 113 -496
rect 104 -503 113 -499
rect 110 -507 113 -503
rect 135 -506 138 -496
rect 155 -506 159 -497
rect 201 -506 205 -423
rect 259 -436 263 -395
rect 864 -422 868 -365
rect 882 -367 892 -365
rect 882 -368 904 -367
rect 889 -370 904 -368
rect 900 -371 904 -370
rect 886 -379 904 -375
rect 885 -387 904 -383
rect 885 -391 889 -387
rect 879 -395 889 -391
rect 893 -395 904 -391
rect 893 -404 897 -395
rect 879 -408 897 -404
rect 900 -411 904 -399
rect 911 -403 915 -343
rect 1042 -351 1079 -347
rect 1083 -348 1086 -343
rect 1083 -351 1093 -348
rect 1042 -355 1046 -351
rect 1039 -359 1046 -355
rect 1061 -359 1068 -355
rect 1042 -363 1046 -359
rect 1042 -367 1051 -363
rect 1042 -379 1046 -367
rect 1064 -371 1068 -359
rect 1061 -375 1068 -371
rect 1042 -383 1051 -379
rect 1042 -395 1046 -383
rect 1064 -387 1068 -375
rect 1075 -383 1079 -351
rect 1089 -354 1093 -351
rect 1275 -354 1318 -350
rect 1238 -361 1247 -357
rect 1097 -383 1101 -374
rect 1136 -365 1231 -361
rect 1075 -387 1090 -383
rect 1097 -387 1107 -383
rect 1061 -391 1068 -387
rect 1097 -390 1101 -387
rect 1042 -399 1051 -395
rect 1064 -402 1068 -391
rect 1124 -395 1128 -382
rect 1136 -395 1140 -365
rect 1227 -384 1231 -369
rect 1238 -373 1241 -361
rect 1275 -365 1279 -354
rect 1303 -361 1306 -357
rect 1267 -369 1279 -365
rect 1275 -373 1279 -369
rect 1184 -388 1231 -384
rect 1147 -395 1156 -391
rect 1124 -399 1140 -395
rect 1089 -402 1093 -400
rect 1064 -403 1093 -402
rect 911 -407 919 -403
rect 1061 -406 1093 -403
rect 1061 -407 1068 -406
rect 903 -416 904 -411
rect 1089 -422 1093 -406
rect 1121 -407 1140 -403
rect 1147 -407 1150 -395
rect 1184 -399 1188 -388
rect 1212 -395 1216 -391
rect 1176 -403 1188 -399
rect 1184 -407 1188 -403
rect 1121 -413 1125 -407
rect 1121 -418 1122 -413
rect 864 -426 1093 -422
rect 110 -511 116 -507
rect 135 -510 148 -506
rect 155 -510 205 -506
rect 210 -439 263 -436
rect 1089 -436 1093 -426
rect 1136 -425 1140 -407
rect 1147 -411 1156 -407
rect 1184 -411 1192 -407
rect 1227 -421 1231 -388
rect 1238 -377 1247 -373
rect 1275 -377 1283 -373
rect 1238 -386 1242 -377
rect 1238 -390 1287 -386
rect 1238 -413 1242 -390
rect 1314 -395 1318 -354
rect 1333 -386 1337 -343
rect 1371 -387 1421 -383
rect 1334 -395 1343 -391
rect 1314 -399 1327 -395
rect 1314 -406 1327 -403
rect 1275 -407 1327 -406
rect 1334 -407 1337 -395
rect 1371 -399 1375 -387
rect 1399 -395 1403 -391
rect 1363 -403 1375 -399
rect 1371 -407 1375 -403
rect 1275 -410 1318 -407
rect 1238 -417 1247 -413
rect 1136 -429 1231 -425
rect 1238 -429 1241 -417
rect 1275 -421 1279 -410
rect 1334 -411 1343 -407
rect 1371 -411 1379 -407
rect 1303 -417 1313 -413
rect 1267 -425 1279 -421
rect 1275 -429 1279 -425
rect 1238 -433 1247 -429
rect 1275 -433 1283 -429
rect 1309 -436 1313 -417
rect 1403 -436 1407 -395
rect 1418 -407 1423 -402
rect 155 -513 159 -510
rect 58 -519 64 -515
rect 126 -519 132 -515
rect 129 -529 132 -519
rect 147 -529 151 -523
rect 210 -529 213 -439
rect 1089 -440 1407 -436
rect 0 -532 213 -529
<< m2contact >>
rect 124 130 129 135
rect 9 78 14 83
rect 30 87 35 92
rect 25 78 30 83
rect 31 63 36 68
rect 25 22 30 27
rect 25 13 30 18
rect 173 118 178 123
rect 45 87 50 92
rect 45 78 50 83
rect 193 118 198 123
rect 46 63 51 68
rect 45 22 50 27
rect 45 13 50 18
rect 162 54 167 59
rect 371 92 376 97
rect 171 41 176 46
rect 177 31 182 36
rect 309 64 314 69
rect 39 4 44 9
rect 177 14 182 19
rect 197 54 202 59
rect 197 41 202 46
rect 212 45 217 50
rect 531 78 536 83
rect 371 49 376 54
rect 331 31 336 36
rect 441 44 446 49
rect 203 9 208 14
rect 342 14 347 19
rect 512 50 517 55
rect 557 49 562 54
rect 628 45 633 50
rect 41 -11 46 -6
rect 127 -7 132 -2
rect 9 -54 14 -49
rect 30 -45 35 -40
rect 25 -54 30 -49
rect 31 -69 36 -64
rect 25 -110 30 -105
rect 25 -119 30 -114
rect 45 -45 50 -40
rect 45 -54 50 -49
rect 177 -21 182 -16
rect 186 -30 191 -25
rect 165 -50 170 -45
rect 318 -22 323 -17
rect 46 -69 51 -64
rect 127 -65 132 -60
rect 306 -50 311 -45
rect 173 -62 178 -57
rect 319 -62 324 -57
rect 625 -18 630 -13
rect 596 -23 601 -18
rect 447 -56 452 -51
rect 583 -50 588 -45
rect 438 -62 443 -57
rect 151 -77 156 -72
rect 183 -76 188 -71
rect 306 -76 311 -71
rect 439 -76 444 -71
rect 448 -76 453 -71
rect 45 -110 50 -105
rect 45 -119 50 -114
rect 173 -84 178 -79
rect 180 -96 185 -91
rect 541 -92 546 -87
rect 196 -108 201 -103
rect 39 -128 44 -123
rect 128 -139 133 -134
rect 39 -144 44 -139
rect 9 -186 14 -181
rect 30 -177 35 -172
rect 25 -186 30 -181
rect 31 -201 36 -196
rect 25 -242 30 -237
rect 25 -251 30 -246
rect 334 -116 339 -111
rect 334 -125 339 -120
rect 183 -144 188 -139
rect 421 -121 426 -116
rect 464 -112 469 -107
rect 785 -32 790 -27
rect 625 -61 630 -56
rect 577 -77 582 -72
rect 695 -66 700 -61
rect 456 -132 461 -127
rect 334 -144 339 -139
rect 766 -60 771 -55
rect 811 -61 816 -56
rect 882 -65 887 -60
rect 585 -120 590 -115
rect 538 -132 543 -127
rect 465 -144 470 -139
rect 45 -177 50 -172
rect 45 -186 50 -181
rect 300 -160 306 -153
rect 425 -158 430 -153
rect 456 -158 461 -153
rect 543 -158 548 -153
rect 179 -168 184 -163
rect 165 -182 170 -177
rect 46 -201 51 -196
rect 128 -197 133 -192
rect 479 -166 484 -161
rect 565 -158 570 -153
rect 778 -128 783 -123
rect 742 -161 747 -156
rect 586 -173 591 -168
rect 938 -142 943 -137
rect 778 -171 783 -166
rect 301 -183 306 -178
rect 326 -183 331 -178
rect 479 -183 484 -178
rect 706 -190 711 -185
rect 157 -202 162 -197
rect 172 -201 177 -196
rect 45 -242 50 -237
rect 45 -251 50 -246
rect 192 -210 197 -205
rect 201 -210 206 -205
rect 188 -237 193 -232
rect 39 -260 44 -255
rect 172 -254 177 -249
rect 281 -242 286 -237
rect 326 -217 331 -212
rect 324 -229 330 -223
rect 472 -212 477 -207
rect 324 -249 329 -244
rect 191 -259 196 -254
rect 287 -257 292 -252
rect 460 -224 465 -219
rect 600 -217 605 -212
rect 424 -250 429 -245
rect 332 -258 337 -253
rect 469 -250 474 -245
rect 733 -190 738 -185
rect 751 -187 756 -182
rect 848 -176 853 -171
rect 919 -170 924 -165
rect 964 -171 969 -166
rect 1035 -175 1040 -170
rect 605 -251 610 -246
rect 677 -247 682 -242
rect 127 -271 132 -266
rect 40 -276 45 -271
rect 202 -274 207 -269
rect 261 -274 266 -269
rect 279 -274 284 -269
rect 332 -274 337 -269
rect 9 -318 14 -313
rect 30 -309 35 -304
rect 25 -318 30 -313
rect 31 -333 36 -328
rect 25 -374 30 -369
rect 25 -383 30 -378
rect 187 -280 192 -275
rect 45 -309 50 -304
rect 45 -318 50 -313
rect 178 -314 183 -309
rect 46 -333 51 -328
rect 127 -329 132 -324
rect 45 -374 50 -369
rect 45 -383 50 -378
rect 226 -307 231 -302
rect 205 -325 210 -320
rect 279 -298 284 -293
rect 702 -259 707 -254
rect 702 -277 707 -272
rect 702 -286 707 -281
rect 939 -237 944 -232
rect 986 -237 991 -232
rect 917 -271 922 -266
rect 1099 -251 1104 -246
rect 939 -280 944 -275
rect 722 -291 727 -286
rect 362 -304 367 -299
rect 208 -359 213 -354
rect 318 -349 323 -344
rect 368 -319 373 -314
rect 360 -333 365 -328
rect 318 -358 323 -353
rect 359 -357 364 -352
rect 39 -392 44 -387
rect 126 -404 131 -399
rect 40 -409 45 -404
rect 9 -451 14 -446
rect 30 -442 35 -437
rect 25 -451 30 -446
rect 31 -466 36 -461
rect 25 -507 30 -502
rect 25 -516 30 -511
rect 177 -411 182 -406
rect 45 -442 50 -437
rect 45 -451 50 -446
rect 210 -411 215 -406
rect 371 -367 377 -361
rect 450 -345 455 -340
rect 485 -335 490 -330
rect 483 -347 488 -342
rect 450 -354 455 -349
rect 597 -344 602 -339
rect 633 -337 638 -332
rect 500 -357 505 -352
rect 597 -353 602 -348
rect 773 -338 778 -333
rect 649 -353 654 -348
rect 906 -290 911 -285
rect 1009 -285 1014 -280
rect 1080 -279 1085 -274
rect 1125 -280 1130 -275
rect 1196 -284 1201 -279
rect 986 -339 991 -334
rect 774 -355 779 -350
rect 245 -423 250 -418
rect 180 -447 185 -442
rect 46 -466 51 -461
rect 126 -462 131 -457
rect 45 -507 50 -502
rect 45 -516 50 -511
rect 1146 -348 1151 -343
rect 1107 -388 1112 -383
rect 1306 -362 1311 -357
rect 1146 -391 1151 -386
rect 898 -416 903 -411
rect 1216 -396 1221 -391
rect 1287 -390 1292 -385
rect 1332 -391 1337 -386
rect 1403 -395 1408 -390
rect 1413 -407 1418 -402
rect 39 -525 44 -520
<< metal2 >>
rect 35 87 45 91
rect 14 79 25 83
rect 30 79 45 83
rect 36 64 46 67
rect 125 42 128 130
rect 178 119 193 123
rect 167 54 197 58
rect 309 50 313 64
rect 372 54 375 92
rect 533 71 536 78
rect 533 68 632 71
rect 533 62 536 68
rect 505 59 536 62
rect 125 39 140 42
rect 176 41 197 45
rect 217 46 313 50
rect 505 48 508 59
rect 517 51 557 54
rect 629 50 632 68
rect 446 45 508 48
rect 30 22 45 25
rect 30 15 45 18
rect 41 -6 44 4
rect 137 -3 140 39
rect 182 31 331 35
rect 137 -6 167 -3
rect 35 -45 45 -41
rect 14 -53 25 -49
rect 30 -53 45 -49
rect 128 -60 131 -7
rect 36 -68 46 -65
rect 137 -103 140 -6
rect 164 -25 167 -6
rect 178 -5 181 14
rect 204 -1 207 9
rect 344 -1 347 14
rect 204 -4 321 -1
rect 344 -4 600 -1
rect 178 -8 199 -5
rect 178 -16 181 -8
rect 164 -28 186 -25
rect 170 -49 186 -46
rect 156 -76 169 -73
rect 166 -92 169 -76
rect 174 -79 177 -62
rect 183 -71 186 -49
rect 196 -70 199 -8
rect 318 -17 321 -4
rect 597 -18 600 -4
rect 307 -71 310 -50
rect 320 -80 323 -62
rect 178 -83 323 -80
rect 393 -83 396 -45
rect 440 -71 443 -62
rect 448 -71 451 -56
rect 584 -62 587 -50
rect 626 -56 629 -18
rect 787 -39 790 -32
rect 787 -42 886 -39
rect 787 -48 790 -42
rect 759 -51 790 -48
rect 584 -65 592 -62
rect 589 -72 592 -65
rect 759 -62 762 -51
rect 771 -59 811 -56
rect 883 -60 886 -42
rect 700 -65 762 -62
rect 453 -75 577 -72
rect 335 -86 396 -83
rect 166 -95 180 -92
rect 30 -110 45 -107
rect 137 -106 196 -103
rect 335 -111 338 -86
rect 465 -107 468 -75
rect 589 -75 601 -72
rect 542 -87 589 -84
rect 30 -117 45 -114
rect 293 -116 296 -113
rect 586 -115 589 -87
rect 598 -95 601 -75
rect 598 -98 607 -95
rect 604 -112 607 -98
rect 604 -115 754 -112
rect 41 -139 44 -128
rect 327 -124 334 -121
rect 327 -135 330 -124
rect 303 -138 330 -135
rect 35 -177 45 -173
rect 14 -185 25 -181
rect 30 -185 45 -181
rect 129 -192 132 -139
rect 180 -163 183 -139
rect 300 -153 303 -139
rect 334 -164 337 -144
rect 426 -153 429 -117
rect 457 -153 460 -132
rect 465 -164 468 -144
rect 543 -146 546 -127
rect 529 -149 546 -146
rect 751 -148 754 -115
rect 184 -167 468 -164
rect 529 -162 532 -149
rect 751 -151 757 -148
rect 548 -157 565 -154
rect 754 -159 757 -151
rect 484 -165 532 -162
rect 289 -174 551 -171
rect 289 -178 292 -174
rect 548 -178 551 -174
rect 587 -178 590 -173
rect 170 -181 292 -178
rect 472 -183 479 -180
rect 548 -181 604 -178
rect 302 -192 305 -183
rect 36 -200 46 -197
rect 185 -195 305 -192
rect 162 -201 172 -198
rect 185 -237 188 -195
rect 327 -203 330 -183
rect 319 -206 330 -203
rect 30 -242 45 -239
rect 30 -249 45 -246
rect 41 -271 44 -260
rect 35 -309 45 -305
rect 14 -317 25 -313
rect 30 -317 45 -313
rect 128 -324 131 -271
rect 173 -295 176 -254
rect 193 -266 196 -259
rect 189 -269 196 -266
rect 203 -269 206 -210
rect 262 -209 322 -206
rect 262 -269 265 -209
rect 327 -212 330 -206
rect 472 -207 475 -183
rect 601 -212 604 -181
rect 711 -189 733 -186
rect 317 -226 324 -223
rect 280 -242 281 -239
rect 317 -238 320 -226
rect 743 -221 746 -161
rect 751 -162 757 -159
rect 751 -182 754 -162
rect 779 -166 782 -128
rect 940 -149 943 -142
rect 940 -152 1039 -149
rect 940 -158 943 -152
rect 912 -161 943 -158
rect 912 -172 915 -161
rect 924 -169 964 -166
rect 1036 -170 1039 -152
rect 853 -175 915 -172
rect 743 -224 930 -221
rect 286 -241 320 -238
rect 280 -269 283 -242
rect 292 -256 308 -253
rect 324 -256 327 -249
rect 460 -246 463 -224
rect 429 -249 463 -246
rect 305 -259 327 -256
rect 469 -257 472 -250
rect 682 -246 921 -243
rect 605 -257 608 -251
rect 333 -269 336 -258
rect 469 -260 608 -257
rect 189 -275 192 -269
rect 469 -270 472 -260
rect 699 -262 702 -255
rect 613 -265 702 -262
rect 337 -273 472 -270
rect 494 -271 538 -268
rect 613 -267 616 -265
rect 918 -266 921 -246
rect 595 -270 616 -267
rect 332 -275 336 -274
rect 298 -278 336 -275
rect 535 -275 538 -271
rect 683 -275 702 -272
rect 192 -280 302 -278
rect 187 -281 302 -280
rect 535 -278 686 -275
rect 927 -275 930 -224
rect 940 -275 943 -237
rect 907 -278 930 -275
rect 360 -281 511 -278
rect 508 -282 511 -281
rect 508 -285 702 -282
rect 907 -285 910 -278
rect 170 -298 176 -295
rect 198 -289 303 -286
rect 36 -332 46 -329
rect 170 -334 173 -298
rect 198 -310 201 -289
rect 300 -291 303 -289
rect 183 -313 201 -310
rect 206 -297 279 -294
rect 206 -320 209 -297
rect 300 -294 672 -291
rect 669 -295 672 -294
rect 722 -295 725 -291
rect 669 -298 776 -295
rect 363 -314 366 -304
rect 363 -317 368 -314
rect 598 -328 636 -325
rect 355 -333 360 -330
rect 170 -337 199 -334
rect 196 -355 199 -337
rect 355 -345 358 -333
rect 451 -334 485 -331
rect 451 -340 454 -334
rect 598 -339 601 -328
rect 633 -332 636 -328
rect 773 -333 776 -298
rect 987 -334 990 -237
rect 1101 -258 1104 -251
rect 1101 -261 1200 -258
rect 1101 -267 1104 -261
rect 1073 -270 1104 -267
rect 1073 -281 1076 -270
rect 1085 -278 1125 -275
rect 1197 -279 1200 -261
rect 1014 -284 1076 -281
rect 323 -348 358 -345
rect 196 -358 208 -355
rect 323 -356 359 -353
rect 483 -350 486 -347
rect 455 -353 486 -350
rect 602 -353 649 -350
rect 501 -365 504 -357
rect 775 -365 778 -355
rect 30 -374 45 -371
rect 371 -377 374 -367
rect 501 -368 778 -365
rect 501 -377 504 -368
rect 30 -381 45 -378
rect 371 -380 504 -377
rect 41 -404 44 -392
rect 371 -398 374 -380
rect 1147 -386 1150 -348
rect 1308 -369 1311 -362
rect 1308 -372 1407 -369
rect 1308 -378 1311 -372
rect 1280 -381 1311 -378
rect 273 -401 331 -398
rect 336 -401 374 -398
rect 35 -442 45 -438
rect 14 -450 25 -446
rect 30 -450 45 -446
rect 127 -457 130 -404
rect 182 -410 210 -407
rect 273 -419 276 -401
rect 250 -422 276 -419
rect 280 -415 869 -412
rect 886 -415 898 -412
rect 280 -429 283 -415
rect 866 -418 889 -415
rect 181 -432 283 -429
rect 181 -442 184 -432
rect 185 -446 186 -443
rect 1108 -445 1111 -388
rect 1280 -392 1283 -381
rect 1292 -389 1332 -386
rect 1404 -390 1407 -372
rect 1221 -395 1283 -392
rect 1413 -445 1416 -407
rect 1108 -448 1416 -445
rect 36 -465 46 -462
rect 30 -507 45 -504
rect 30 -514 45 -511
<< m3contact >>
rect 195 -75 200 -70
rect 293 -121 298 -116
rect 313 -251 319 -245
rect 489 -272 494 -267
rect 590 -271 595 -266
rect 355 -282 360 -277
<< metal3 >>
rect 196 -96 199 -75
rect 190 -99 199 -96
rect 190 -116 193 -99
rect 190 -156 193 -121
rect 184 -159 193 -156
rect 184 -217 187 -159
rect 293 -171 296 -121
rect 321 -130 329 -127
rect 326 -159 329 -130
rect 326 -162 564 -159
rect 561 -164 564 -162
rect 561 -167 568 -164
rect 193 -174 296 -171
rect 193 -205 196 -174
rect 184 -220 192 -217
rect 184 -303 187 -220
rect 314 -278 318 -251
rect 459 -268 462 -258
rect 459 -271 489 -268
rect 314 -282 355 -278
rect 555 -293 558 -228
rect 590 -266 593 -239
rect 498 -296 558 -293
rect 184 -306 226 -303
rect 498 -313 501 -296
rect 678 -300 681 -230
rect 906 -266 1129 -263
rect 643 -303 681 -300
rect 643 -316 646 -303
rect 330 -352 368 -349
rect 330 -364 333 -352
rect 323 -367 333 -364
rect 332 -418 335 -403
rect 355 -405 358 -385
rect 473 -391 476 -364
rect 630 -380 633 -346
rect 766 -372 769 -347
rect 871 -370 877 -367
rect 871 -372 874 -370
rect 766 -375 874 -372
rect 878 -380 881 -375
rect 1126 -377 1129 -266
rect 630 -383 881 -380
rect 473 -394 874 -391
rect 355 -408 874 -405
rect 332 -421 855 -418
rect 852 -428 855 -421
rect 1122 -428 1125 -418
rect 852 -431 1125 -428
<< labels >>
rlabel metal1 -1 119 2 122 4 VDD
rlabel metal1 161 83 165 87 7 G0
rlabel metal1 161 19 165 23 7 P0
rlabel metal1 161 -49 165 -45 7 G1
rlabel metal1 161 -113 165 -109 7 P1
rlabel metal1 161 -181 165 -177 7 G2
rlabel metal1 161 -245 165 -241 7 P2
rlabel metal1 161 -377 165 -373 7 P3
rlabel metal1 161 -510 165 -506 7 P4
rlabel metal1 0 -532 3 -529 2 GND
rlabel metal1 0 88 9 97 3 A0
rlabel metal1 0 74 9 83 3 B0
rlabel metal1 0 -44 9 -35 3 A1
rlabel metal1 0 -58 9 -49 3 B1
rlabel metal1 0 -176 9 -167 3 A2
rlabel metal1 0 -190 9 -181 3 B2
rlabel metal1 0 -308 9 -299 3 A3
rlabel metal1 0 -322 9 -313 3 B3
rlabel metal1 0 -441 9 -432 3 A4
rlabel metal1 0 -455 9 -446 3 B4
rlabel metal1 -1 135 8 144 4 Cin
rlabel metal1 323 19 327 23 7 C1
rlabel metal1 642 53 646 57 7 S0
rlabel metal1 579 -49 583 -45 1 C2
rlabel metal1 896 -57 900 -53 7 S1
rlabel metal1 740 -160 744 -156 1 C3
rlabel metal1 1049 -167 1053 -163 7 S2
rlabel metal1 160 -313 164 -309 1 G3
rlabel metal1 897 -266 901 -262 1 C4
rlabel metal1 1210 -276 1214 -272 7 S3
rlabel metal1 1103 -387 1107 -383 1 C5
rlabel metal1 161 -446 165 -442 7 G4
rlabel metal1 1417 -387 1421 -383 7 S4
rlabel metal1 1418 -407 1423 -402 7 Cout
<< end >>
