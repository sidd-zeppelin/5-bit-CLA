* NGSPICE file created from OR6.ext - technology: scmos

.global Vdd Gnd 


* Top level circuit OR6

M1000 a_19_47# C GND Gnd cmosn w=0.9u l=0.18u
+  ad=1.458p pd=8.64u as=2.187p ps=13.86u
M1001 OUT a_19_47# GND Gnd cmosn w=0.9u l=0.18u
+  ad=0.405p pd=2.7u as=0p ps=0u
M1002 a_19_47# A GND Gnd cmosn w=0.9u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1003 GND F a_19_47# Gnd cmosn w=0.9u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1004 OUT a_19_47# VDD w_183_27# cmosp w=1.8u l=0.18u
+  ad=0.81p pd=4.5u as=5.67p ps=27u
M1005 a_19_7# A VDD w_13_n6# cmosp w=10.8u l=0.18u
+  ad=5.832p pd=22.68u as=0p ps=0u
M1006 a_19_31# D a_19_23# w_13_n6# cmosp w=10.8u l=0.18u
+  ad=5.832p pd=22.68u as=5.832p ps=22.68u
M1007 a_19_15# B a_19_7# w_13_n6# cmosp w=10.8u l=0.18u
+  ad=5.832p pd=22.68u as=0p ps=0u
M1008 GND D a_19_47# Gnd cmosn w=0.9u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1009 a_19_39# E a_19_31# w_13_n6# cmosp w=10.8u l=0.18u
+  ad=5.832p pd=22.68u as=0p ps=0u
M1010 GND B a_19_47# Gnd cmosn w=0.9u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_19_23# C a_19_15# w_13_n6# cmosp w=10.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_19_47# E GND Gnd cmosn w=0.9u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_19_47# F a_19_39# w_13_n6# cmosp w=10.8u l=0.18u
+  ad=4.86p pd=22.5u as=0p ps=0u
.end

