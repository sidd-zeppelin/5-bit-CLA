magic
tech scmos
timestamp 1764767778
<< nwell >>
rect 5 -9 97 39
<< polysilicon >>
rect 2 26 11 28
rect 91 26 103 28
rect 113 26 116 28
rect 2 18 11 20
rect 91 18 103 20
rect 113 18 116 20
rect 2 10 11 12
rect 91 10 103 12
rect 113 10 116 12
rect 2 2 11 4
rect 91 2 103 4
rect 113 2 116 4
<< ndiffusion >>
rect 103 28 113 29
rect 103 25 113 26
rect 103 20 113 21
rect 103 17 113 18
rect 103 12 113 13
rect 103 9 113 10
rect 103 4 113 5
rect 103 1 113 2
<< pdiffusion >>
rect 11 28 91 29
rect 11 25 91 26
rect 11 20 91 21
rect 11 17 91 18
rect 11 12 91 13
rect 11 9 91 10
rect 11 4 91 5
rect 11 1 91 2
<< metal1 >>
rect -6 25 -2 29
rect -6 17 -2 21
rect -6 9 -2 13
rect -6 1 -2 5
rect 5 1 8 39
rect 96 36 122 39
rect 96 33 99 36
rect 91 29 99 33
rect 113 29 119 33
rect 95 25 99 29
rect 95 21 103 25
rect 95 9 99 21
rect 116 17 119 29
rect 113 13 119 17
rect 95 5 103 9
rect 116 1 119 13
rect 5 -3 11 1
rect 113 -3 119 1
rect 5 -9 8 -3
<< ntransistor >>
rect 103 26 113 28
rect 103 18 113 20
rect 103 10 113 12
rect 103 2 113 4
<< ptransistor >>
rect 11 26 91 28
rect 11 18 91 20
rect 11 10 91 12
rect 11 2 91 4
<< polycontact >>
rect -2 25 2 29
rect -2 17 2 21
rect -2 9 2 13
rect -2 1 2 5
<< ndcontact >>
rect 103 29 113 33
rect 103 21 113 25
rect 103 13 113 17
rect 103 5 113 9
rect 103 -3 113 1
<< pdcontact >>
rect 11 29 91 33
rect 11 21 91 25
rect 11 13 91 17
rect 11 5 91 9
rect 11 -3 91 1
<< labels >>
rlabel metal1 -6 1 -2 5 3 A
rlabel metal1 -6 9 -2 13 3 B
rlabel metal1 -6 17 -2 21 3 C
rlabel metal1 -6 25 -2 29 3 D
rlabel metal1 5 -9 8 39 7 VDD
rlabel metal1 116 -3 119 33 7 GND
rlabel metal1 119 36 122 39 6 OUT
<< end >>
