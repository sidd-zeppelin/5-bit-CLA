* NGSPICE file created from master_slave_D_FF.ext - technology: scmos

.global Vdd Gnd 


* Top level circuit master_slave_D_FF

M1000 GND a_n22_n1# a_120_17# Gnd cmosn w=1.8u l=0.18u
+  ad=8.1p pd=46.8u as=0.972p ps=4.68u
M1001 GND a_n111_n64# a_14_n48# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1002 a_341_n48# a_267_n64# a_305_n48# Gnd cmosn w=1.8u l=0.18u
+  ad=0.972p pd=4.68u as=0.81p ps=4.5u
M1003 a_n111_n64# CLK VDD w_n124_n46# cmosp w=1.8u l=0.18u
+  ad=0.81p pd=4.5u as=16.2p ps=90u
M1004 a_217_n64# a_n111_n64# VDD w_204_n46# cmosp w=1.8u l=0.18u
+  ad=0.81p pd=4.5u as=0p ps=0u
M1005 a_n60_n64# D_in GND Gnd cmosn w=0.9u l=0.18u
+  ad=0.405p pd=2.7u as=0p ps=0u
M1006 a_68_14# a_n22_n48# VDD w_78_n61# cmosp w=1.8u l=0.18u
+  ad=0.972p pd=4.68u as=0p ps=0u
M1007 VDD a_305_n1# Q w_405_4# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1008 a_68_n43# a_68_14# VDD w_78_4# cmosp w=1.8u l=0.18u
+  ad=0.972p pd=4.68u as=0p ps=0u
M1009 VDD a_n111_n64# a_n22_n48# w_n28_n61# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1010 VDD a_68_n43# a_305_n1# w_299_n14# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1011 a_447_n48# a_305_n48# a_395_14# Gnd cmosn w=1.8u l=0.18u
+  ad=0.972p pd=4.68u as=0.81p ps=4.5u
M1012 a_n111_n64# CLK GND Gnd cmosn w=0.9u l=0.18u
+  ad=0.405p pd=2.7u as=0p ps=0u
M1013 VDD D_in a_n22_n1# w_n28_n14# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1014 a_305_n1# a_217_n64# VDD w_299_n14# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1015 VDD a_217_n64# a_305_n48# w_299_n61# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1016 a_120_n48# a_n22_n48# a_68_14# Gnd cmosn w=1.8u l=0.18u
+  ad=0.972p pd=4.68u as=0.81p ps=4.5u
M1017 a_217_n64# a_n111_n64# GND Gnd cmosn w=0.9u l=0.18u
+  ad=0.405p pd=2.7u as=0p ps=0u
M1018 a_395_14# a_305_n48# VDD w_405_n61# cmosp w=1.8u l=0.18u
+  ad=0.972p pd=4.68u as=0p ps=0u
M1019 GND a_68_n43# a_341_n1# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1020 a_14_n1# a_n111_n64# a_n22_n1# Gnd cmosn w=1.8u l=0.18u
+  ad=0.972p pd=4.68u as=0.81p ps=4.5u
M1021 GND a_217_n64# a_341_n48# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1022 VDD a_n22_n1# a_68_n43# w_78_4# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1023 a_447_17# a_395_14# Q Gnd cmosn w=1.8u l=0.18u
+  ad=0.972p pd=4.68u as=0.81p ps=4.5u
M1024 a_14_n48# a_n60_n64# a_n22_n48# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.81p ps=4.5u
M1025 VDD a_68_n43# a_68_14# w_78_n61# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1026 a_267_n64# a_68_n43# VDD w_254_n46# cmosp w=1.8u l=0.18u
+  ad=0.81p pd=4.5u as=0p ps=0u
M1027 a_120_17# a_68_14# a_68_n43# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.81p ps=4.5u
M1028 GND Q a_447_n48# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1029 a_n22_n48# a_n60_n64# VDD w_n28_n61# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1030 GND a_68_n43# a_120_n48# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1031 VDD Q a_395_14# w_405_n61# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1032 GND a_305_n1# a_447_17# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1033 GND D_in a_14_n1# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1034 a_n60_n64# D_in VDD w_n73_n46# cmosp w=1.8u l=0.18u
+  ad=0.81p pd=4.5u as=0p ps=0u
M1035 a_305_n48# a_267_n64# VDD w_299_n61# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1036 a_267_n64# a_68_n43# GND Gnd cmosn w=0.9u l=0.18u
+  ad=0.405p pd=2.7u as=0p ps=0u
M1037 Q a_395_14# VDD w_405_4# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1038 a_n22_n1# a_n111_n64# VDD w_n28_n14# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1039 a_341_n1# a_217_n64# a_305_n1# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.81p ps=4.5u
.end

