magic
tech scmos
timestamp 1764685615
<< nwell >>
rect -27 107 5 131
rect 55 107 87 131
rect -6 28 42 80
<< ntransistor >>
rect -47 118 -37 120
rect 35 118 45 120
rect 5 0 7 20
rect 13 0 15 20
rect 21 0 23 20
rect 29 0 31 20
<< ptransistor >>
rect -21 118 -1 120
rect 61 118 81 120
rect 5 34 7 74
rect 13 34 15 74
rect 21 34 23 74
rect 29 34 31 74
<< ndiffusion >>
rect -47 120 -37 121
rect 35 120 45 121
rect -47 117 -37 118
rect 35 117 45 118
rect 4 0 5 20
rect 7 0 8 20
rect 12 0 13 20
rect 15 0 16 20
rect 20 0 21 20
rect 23 0 24 20
rect 28 0 29 20
rect 31 0 33 20
<< pdiffusion >>
rect -21 120 -1 121
rect 61 120 81 121
rect -21 117 -1 118
rect 61 117 81 118
rect 4 34 5 74
rect 7 34 8 74
rect 12 34 13 74
rect 15 34 16 74
rect 20 34 21 74
rect 23 34 24 74
rect 28 34 29 74
rect 31 34 32 74
<< ndcontact >>
rect -47 121 -37 125
rect 35 121 45 125
rect -47 113 -37 117
rect 35 113 45 117
rect 0 0 4 20
rect 8 0 12 20
rect 16 0 20 20
rect 24 0 28 20
rect 33 0 37 20
<< pdcontact >>
rect -21 121 -1 125
rect 61 121 81 125
rect -21 113 -1 117
rect 61 113 81 117
rect 0 34 4 74
rect 8 34 12 74
rect 16 34 20 74
rect 24 34 28 74
rect 32 34 36 74
<< polysilicon >>
rect -50 118 -47 120
rect -37 118 -21 120
rect -1 118 2 120
rect 32 118 35 120
rect 45 118 61 120
rect 81 118 84 120
rect 5 74 7 84
rect 13 74 15 84
rect 21 74 23 84
rect 29 74 31 84
rect 5 20 7 34
rect 13 20 15 34
rect 21 20 23 34
rect 29 20 31 34
rect 5 -3 7 0
rect 13 -3 15 0
rect 21 -3 23 0
rect 29 -3 31 0
<< polycontact >>
rect -34 120 -30 124
rect 48 120 52 124
rect 4 84 8 88
rect 12 84 16 88
rect 20 84 24 88
rect 28 84 32 88
<< metal1 >>
rect -34 138 16 142
rect -53 121 -47 125
rect -34 124 -30 138
rect 2 125 5 131
rect -53 113 -50 121
rect -1 121 5 125
rect -37 113 -21 117
rect -34 96 -30 113
rect 2 107 5 121
rect -34 92 8 96
rect 4 88 8 92
rect 12 88 16 138
rect 48 138 94 142
rect 29 121 35 125
rect 48 124 52 138
rect 84 125 87 131
rect 29 113 32 121
rect 81 121 87 125
rect 45 113 61 117
rect 48 96 52 113
rect 84 107 87 121
rect 20 92 52 96
rect 20 88 24 92
rect 90 88 94 138
rect 32 84 94 88
rect 0 77 36 81
rect 0 74 4 77
rect 16 74 20 77
rect 32 74 36 77
rect 8 30 12 34
rect 24 30 28 34
rect -6 26 12 30
rect 16 26 28 30
rect 16 20 20 26
rect 0 -3 4 0
rect 33 -3 37 0
rect -6 -7 37 -3
<< labels >>
rlabel metal1 -6 26 -2 30 3 VDD
rlabel metal1 -6 -7 -2 -3 2 GND
rlabel metal1 -34 127 -30 131 5 A
rlabel metal1 -34 107 -30 111 1 OUT
rlabel metal1 -53 113 -50 125 3 GND
rlabel metal1 2 107 5 131 7 VDD
rlabel metal1 48 127 52 131 5 A
rlabel metal1 48 107 52 111 1 OUT
rlabel metal1 29 113 32 125 3 GND
rlabel metal1 84 107 87 131 7 VDD
<< end >>
