* SPICE3 file created from OR2.ext - technology: scmos

.option scale=0.09u

M1000 OUT a_17_21# GND Gnd cmosn w=10 l=2
+  ad=50 pd=30 as=100 ps=60
M1001 a_17_21# A GND Gnd cmosn w=10 l=2
+  ad=60 pd=32 as=0 ps=0
M1002 a_17_21# B a_17_13# w_11_0# cmosp w=40 l=2
+  ad=200 pd=90 as=240 ps=92
M1003 OUT a_17_21# VDD w_94_22# cmosp w=20 l=2
+  ad=100 pd=50 as=300 ps=140
M1004 a_69_21# B a_17_21# Gnd cmosn w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1005 a_17_13# A VDD w_11_0# cmosp w=40 l=2
+  ad=0 pd=0 as=0 ps=0
