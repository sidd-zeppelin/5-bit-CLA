magic
tech scmos
timestamp 1763737113
<< nwell >>
rect -27 -29 5 3
rect 46 -8 70 24
<< ntransistor >>
rect 12 -10 32 -8
rect 12 -18 32 -16
rect 57 -28 59 -18
<< ptransistor >>
rect 57 -2 59 18
rect -21 -10 -1 -8
rect -21 -18 -1 -16
<< ndiffusion >>
rect 12 -8 32 -7
rect 12 -11 32 -10
rect 12 -16 32 -15
rect 12 -19 32 -18
rect 56 -28 57 -18
rect 59 -28 60 -18
<< pdiffusion >>
rect 56 -2 57 18
rect 59 -2 60 18
rect -21 -8 -1 -7
rect -21 -11 -1 -10
rect -21 -16 -1 -15
rect -21 -19 -1 -18
<< ndcontact >>
rect 12 -7 32 -3
rect 12 -15 32 -11
rect 12 -23 32 -19
rect 52 -28 56 -18
rect 60 -28 64 -18
<< pdcontact >>
rect 52 -2 56 18
rect 60 -2 64 18
rect -21 -7 -1 -3
rect -21 -15 -1 -11
rect -21 -23 -1 -19
<< polysilicon >>
rect 57 18 59 21
rect -30 -10 -21 -8
rect -1 -10 12 -8
rect 32 -10 35 -8
rect -30 -18 -21 -16
rect -1 -18 12 -16
rect 32 -18 35 -16
rect 57 -18 59 -2
rect 57 -31 59 -28
<< polycontact >>
rect -34 -11 -30 -7
rect -34 -19 -30 -15
rect 53 -15 57 -11
<< metal1 >>
rect -38 21 56 24
rect -27 -3 -24 21
rect 52 18 56 21
rect 5 0 45 4
rect 5 -3 9 0
rect -27 -7 -21 -3
rect 5 -7 12 -3
rect -38 -11 -34 -7
rect -38 -19 -34 -15
rect -27 -19 -24 -7
rect 5 -11 9 -7
rect 41 -11 45 0
rect 60 -11 64 -2
rect -1 -15 9 -11
rect 41 -15 53 -11
rect 60 -15 70 -11
rect 60 -18 64 -15
rect -27 -23 -21 -19
rect 32 -23 38 -19
rect 35 -31 38 -23
rect 52 -31 56 -28
rect -38 -34 56 -31
<< labels >>
rlabel metal1 -27 -23 -24 -3 3 VDD
rlabel metal1 -38 -19 -34 -15 3 A
rlabel metal1 -38 -11 -34 -7 3 B
rlabel metal1 66 -15 70 -11 7 OUT
rlabel metal1 -38 21 -33 24 4 VDD
rlabel metal1 -38 -34 -33 -31 2 GND
<< end >>
