magic
tech scmos
timestamp 1764589602
<< nwell >>
rect 13 -6 145 58
rect 183 27 207 59
<< ntransistor >>
rect 151 45 161 47
rect 151 37 161 39
rect 151 29 161 31
rect 151 21 161 23
rect 151 13 161 15
rect 194 7 196 17
rect 151 5 161 7
<< ptransistor >>
rect 19 45 139 47
rect 19 37 139 39
rect 194 33 196 53
rect 19 29 139 31
rect 19 21 139 23
rect 19 13 139 15
rect 19 5 139 7
<< ndiffusion >>
rect 151 47 161 48
rect 151 44 161 45
rect 151 39 161 40
rect 151 36 161 37
rect 151 31 161 32
rect 151 28 161 29
rect 151 23 161 24
rect 151 20 161 21
rect 151 15 161 16
rect 151 12 161 13
rect 151 7 161 8
rect 193 7 194 17
rect 196 7 197 17
rect 151 4 161 5
<< pdiffusion >>
rect 19 47 139 48
rect 19 44 139 45
rect 19 39 139 40
rect 19 36 139 37
rect 19 31 139 32
rect 193 33 194 53
rect 196 33 197 53
rect 19 28 139 29
rect 19 23 139 24
rect 19 20 139 21
rect 19 15 139 16
rect 19 12 139 13
rect 19 7 139 8
rect 19 4 139 5
<< ndcontact >>
rect 151 48 161 52
rect 151 40 161 44
rect 151 32 161 36
rect 151 24 161 28
rect 151 16 161 20
rect 151 8 161 12
rect 189 7 193 17
rect 197 7 201 17
rect 151 0 161 4
<< pdcontact >>
rect 19 48 139 52
rect 19 40 139 44
rect 19 32 139 36
rect 189 33 193 53
rect 197 33 201 53
rect 19 24 139 28
rect 19 16 139 20
rect 19 8 139 12
rect 19 0 139 4
<< polysilicon >>
rect 194 53 196 56
rect 8 45 19 47
rect 139 45 151 47
rect 161 45 164 47
rect 8 37 19 39
rect 139 37 151 39
rect 161 37 164 39
rect 8 29 19 31
rect 139 29 151 31
rect 161 29 164 31
rect 8 21 19 23
rect 139 21 151 23
rect 161 21 164 23
rect 194 17 196 33
rect 8 13 19 15
rect 139 13 151 15
rect 161 13 164 15
rect 8 5 19 7
rect 139 5 151 7
rect 161 5 164 7
rect 194 4 196 7
<< polycontact >>
rect 4 44 8 48
rect 4 36 8 40
rect 4 28 8 32
rect 4 20 8 24
rect 4 12 8 16
rect 190 20 194 24
rect 4 4 8 8
<< metal1 >>
rect 11 64 186 68
rect 0 44 4 48
rect 0 36 4 40
rect 0 28 4 32
rect 0 20 4 24
rect 0 12 4 16
rect 0 4 4 8
rect 11 4 15 64
rect 142 56 179 60
rect 183 59 186 64
rect 183 56 193 59
rect 142 52 146 56
rect 139 48 146 52
rect 161 48 168 52
rect 142 44 146 48
rect 142 40 151 44
rect 142 28 146 40
rect 164 36 168 48
rect 161 32 168 36
rect 142 24 151 28
rect 142 12 146 24
rect 164 20 168 32
rect 175 24 179 56
rect 189 53 193 56
rect 197 24 201 33
rect 175 20 190 24
rect 197 20 207 24
rect 161 16 168 20
rect 197 17 201 20
rect 142 8 151 12
rect 164 5 168 16
rect 189 5 193 7
rect 164 4 193 5
rect 11 0 19 4
rect 161 1 193 4
rect 161 0 168 1
<< labels >>
rlabel metal1 0 4 4 8 3 A
rlabel metal1 0 12 4 16 3 B
rlabel metal1 0 20 4 24 3 C
rlabel metal1 0 28 4 32 3 D
rlabel metal1 0 36 4 40 3 E
rlabel metal1 0 44 4 48 3 F
rlabel metal1 203 20 207 24 7 OUT
rlabel metal1 189 1 193 5 1 GND
rlabel metal1 11 0 15 4 1 VDD
<< end >>
