magic
tech scmos
timestamp 1763729104
<< nwell >>
rect 5 -11 37 21
<< ntransistor >>
rect 44 8 64 10
rect 44 0 64 2
<< ptransistor >>
rect 11 8 31 10
rect 11 0 31 2
<< ndiffusion >>
rect 44 10 64 11
rect 44 7 64 8
rect 44 2 64 3
rect 44 -1 64 0
<< pdiffusion >>
rect 11 10 31 11
rect 11 7 31 8
rect 11 2 31 3
rect 11 -1 31 0
<< ndcontact >>
rect 44 11 64 15
rect 44 3 64 7
rect 44 -5 64 -1
<< pdcontact >>
rect 11 11 31 15
rect 11 3 31 7
rect 11 -5 31 -1
<< polysilicon >>
rect 2 8 11 10
rect 31 8 44 10
rect 64 8 67 10
rect 2 0 11 2
rect 31 0 44 2
rect 64 0 67 2
<< polycontact >>
rect -2 7 2 11
rect -2 -1 2 3
<< metal1 >>
rect 37 18 74 22
rect 37 15 41 18
rect 5 11 11 15
rect 37 11 44 15
rect -6 7 -2 11
rect -6 -1 -2 3
rect 5 -1 8 11
rect 37 7 41 11
rect 31 3 41 7
rect 67 -1 70 15
rect 5 -5 11 -1
rect 64 -5 70 -1
<< labels >>
rlabel metal1 5 -5 8 15 3 VDD
rlabel metal1 -6 -1 -2 3 3 A
rlabel metal1 -6 7 -2 11 3 B
rlabel metal1 67 -5 70 15 7 GND
rlabel metal1 70 18 74 22 6 OUT
<< end >>
