magic
tech scmos
timestamp 1763746981
<< nwell >>
rect -6 31 50 63
<< ntransistor >>
rect 5 0 7 25
rect 13 0 15 25
rect 21 0 23 25
rect 29 0 31 25
rect 37 0 39 25
<< ptransistor >>
rect 5 37 7 57
rect 13 37 15 57
rect 21 37 23 57
rect 29 37 31 57
rect 37 37 39 57
<< ndiffusion >>
rect 4 0 5 25
rect 7 0 8 25
rect 12 0 13 25
rect 15 0 16 25
rect 20 0 21 25
rect 23 0 24 25
rect 28 0 29 25
rect 31 0 32 25
rect 36 0 37 25
rect 39 0 40 25
<< pdiffusion >>
rect 4 37 5 57
rect 7 37 8 57
rect 12 37 13 57
rect 15 37 16 57
rect 20 37 21 57
rect 23 37 24 57
rect 28 37 29 57
rect 31 37 32 57
rect 36 37 37 57
rect 39 37 40 57
<< ndcontact >>
rect 0 0 4 25
rect 8 0 12 25
rect 16 0 20 25
rect 24 0 28 25
rect 32 0 36 25
rect 40 0 44 25
<< pdcontact >>
rect 0 37 4 57
rect 8 37 12 57
rect 16 37 20 57
rect 24 37 28 57
rect 32 37 36 57
rect 40 37 44 57
<< polysilicon >>
rect 5 57 7 66
rect 13 57 15 66
rect 21 57 23 66
rect 29 57 31 66
rect 37 57 39 66
rect 5 25 7 37
rect 13 25 15 37
rect 21 25 23 37
rect 29 25 31 37
rect 37 25 39 37
rect 5 -3 7 0
rect 13 -3 15 0
rect 21 -3 23 0
rect 29 -3 31 0
rect 37 -3 39 0
<< polycontact >>
rect 4 66 8 70
rect 12 66 16 70
rect 20 66 24 70
rect 28 66 32 70
rect 36 66 40 70
<< metal1 >>
rect 4 70 8 74
rect 12 70 16 74
rect 20 70 24 74
rect 28 70 32 74
rect 36 70 40 74
rect -6 60 50 63
rect 0 57 4 60
rect 16 57 20 60
rect 32 57 36 60
rect 8 32 12 37
rect 24 32 28 37
rect 40 32 44 37
rect 8 31 44 32
rect 8 28 50 31
rect 40 25 44 28
rect 0 -3 4 0
rect 0 -6 44 -3
rect 47 -9 50 28
<< labels >>
rlabel metal1 0 -6 44 -3 1 GND
rlabel metal1 -6 60 50 63 5 VDD
rlabel metal1 4 70 8 74 5 A
rlabel metal1 12 70 16 74 5 B
rlabel metal1 20 70 24 74 5 C
rlabel metal1 28 70 32 74 5 D
rlabel metal1 36 70 40 74 5 E
rlabel metal1 47 -9 50 -6 8 OUT
<< end >>
