magic
tech scmos
timestamp 1764748415
<< nwell >>
rect 408 207 440 239
rect 317 173 349 205
rect 408 151 440 183
rect 504 173 536 205
rect 157 119 189 151
rect 66 85 98 117
rect 157 63 189 95
rect 253 85 285 117
rect 360 66 392 98
rect 433 87 457 119
rect 478 65 530 97
rect 561 87 585 119
rect 51 5 83 37
rect 124 26 148 58
rect 283 -20 315 12
rect 356 1 380 33
rect 407 -25 479 15
rect 509 -6 533 26
rect 156 -61 188 -29
rect 65 -95 97 -63
rect 156 -117 188 -85
rect 252 -95 284 -63
rect 366 -110 398 -70
rect 448 -92 472 -60
rect 50 -175 82 -143
rect 123 -154 147 -122
rect 647 -148 679 -116
rect 288 -188 320 -156
rect 556 -182 588 -150
rect 197 -222 229 -190
rect 288 -244 320 -212
rect 384 -222 416 -190
rect 647 -204 679 -172
rect 743 -182 775 -150
rect 156 -315 188 -283
rect 540 -286 572 -254
rect 613 -265 637 -233
rect 65 -349 97 -317
rect 156 -371 188 -339
rect 252 -349 284 -317
rect 371 -353 403 -305
rect 463 -330 487 -298
rect 540 -347 572 -307
rect 622 -329 646 -297
rect 687 -339 779 -291
rect 810 -318 834 -286
rect 50 -429 82 -397
rect 123 -408 147 -376
rect 717 -407 749 -375
rect 790 -386 814 -354
rect 157 -497 189 -465
rect 299 -474 331 -418
rect 377 -442 401 -410
rect 435 -464 467 -416
rect 527 -441 551 -409
rect 581 -459 613 -419
rect 663 -441 687 -409
rect 727 -495 839 -439
rect 868 -462 892 -430
rect 66 -531 98 -499
rect 157 -553 189 -521
rect 253 -531 285 -499
rect 51 -611 83 -579
rect 124 -590 148 -558
rect 480 -566 512 -534
rect 389 -600 421 -568
rect 480 -622 512 -590
rect 576 -600 608 -568
rect 698 -627 730 -587
rect 780 -609 804 -577
rect 844 -607 876 -575
rect 917 -586 941 -554
rect 1105 -569 1137 -537
rect 1014 -603 1046 -571
rect 1105 -625 1137 -593
rect 1201 -603 1233 -571
rect 158 -680 190 -648
rect 67 -714 99 -682
rect 158 -736 190 -704
rect 254 -714 286 -682
rect 380 -722 403 -658
rect 462 -689 486 -657
rect 517 -712 549 -656
rect 595 -680 619 -648
rect 645 -712 677 -664
rect 737 -689 761 -657
rect 856 -724 988 -660
rect 1026 -691 1050 -659
rect 52 -794 84 -762
rect 125 -773 149 -741
<< ntransistor >>
rect 450 226 470 228
rect 450 218 470 220
rect 359 192 379 194
rect 546 192 566 194
rect 359 184 379 186
rect 546 184 566 186
rect 450 170 470 172
rect 450 162 470 164
rect 199 138 219 140
rect 199 130 219 132
rect 108 104 128 106
rect 295 104 315 106
rect 108 96 128 98
rect 295 96 315 98
rect 399 85 419 87
rect 199 82 219 84
rect 399 77 419 79
rect 536 84 546 86
rect 199 74 219 76
rect 444 67 446 77
rect 536 76 546 78
rect 572 67 574 77
rect 90 24 110 26
rect 90 16 110 18
rect 135 6 137 16
rect 322 -1 342 1
rect 322 -9 342 -7
rect 485 2 495 4
rect 485 -6 495 -4
rect 367 -19 369 -9
rect 485 -14 495 -12
rect 520 -26 522 -16
rect 198 -42 218 -40
rect 198 -50 218 -48
rect 107 -76 127 -74
rect 294 -76 314 -74
rect 107 -84 127 -82
rect 294 -84 314 -82
rect 404 -83 434 -81
rect 404 -91 434 -89
rect 198 -98 218 -96
rect 404 -99 434 -97
rect 198 -106 218 -104
rect 459 -112 461 -102
rect 689 -129 709 -127
rect 689 -137 709 -135
rect 89 -156 109 -154
rect 89 -164 109 -162
rect 134 -174 136 -164
rect 598 -163 618 -161
rect 330 -169 350 -167
rect 785 -163 805 -161
rect 598 -171 618 -169
rect 330 -177 350 -175
rect 785 -171 805 -169
rect 689 -185 709 -183
rect 689 -193 709 -191
rect 239 -203 259 -201
rect 426 -203 446 -201
rect 239 -211 259 -209
rect 426 -211 446 -209
rect 330 -225 350 -223
rect 330 -233 350 -231
rect 579 -267 599 -265
rect 579 -275 599 -273
rect 624 -285 626 -275
rect 198 -296 218 -294
rect 198 -304 218 -302
rect 409 -318 449 -316
rect 107 -330 127 -328
rect 578 -320 608 -318
rect 409 -326 449 -324
rect 294 -330 314 -328
rect 107 -338 127 -336
rect 409 -334 449 -332
rect 294 -338 314 -336
rect 785 -304 795 -302
rect 785 -312 795 -310
rect 785 -320 795 -318
rect 578 -328 608 -326
rect 578 -336 608 -334
rect 409 -342 449 -340
rect 474 -350 476 -340
rect 785 -328 795 -326
rect 821 -338 823 -328
rect 633 -349 635 -339
rect 198 -352 218 -350
rect 198 -360 218 -358
rect 756 -388 776 -386
rect 756 -396 776 -394
rect 89 -410 109 -408
rect 89 -418 109 -416
rect 801 -406 803 -396
rect 134 -428 136 -418
rect 337 -431 362 -429
rect 473 -429 513 -427
rect 337 -439 362 -437
rect 337 -447 362 -445
rect 619 -432 649 -430
rect 473 -437 513 -435
rect 473 -445 513 -443
rect 337 -455 362 -453
rect 337 -463 362 -461
rect 388 -462 390 -452
rect 619 -440 649 -438
rect 619 -448 649 -446
rect 473 -453 513 -451
rect 538 -461 540 -451
rect 674 -461 676 -451
rect 845 -452 855 -450
rect 845 -460 855 -458
rect 845 -468 855 -466
rect 199 -478 219 -476
rect 845 -476 855 -474
rect 199 -486 219 -484
rect 879 -482 881 -472
rect 845 -484 855 -482
rect 108 -512 128 -510
rect 295 -512 315 -510
rect 108 -520 128 -518
rect 295 -520 315 -518
rect 199 -534 219 -532
rect 199 -542 219 -540
rect 522 -547 542 -545
rect 1147 -550 1167 -548
rect 522 -555 542 -553
rect 1147 -558 1167 -556
rect 431 -581 451 -579
rect 90 -592 110 -590
rect 90 -600 110 -598
rect 618 -581 638 -579
rect 431 -589 451 -587
rect 618 -589 638 -587
rect 135 -610 137 -600
rect 736 -600 766 -598
rect 522 -603 542 -601
rect 883 -588 903 -586
rect 883 -596 903 -594
rect 1056 -584 1076 -582
rect 1243 -584 1263 -582
rect 1056 -592 1076 -590
rect 736 -608 766 -606
rect 522 -611 542 -609
rect 736 -616 766 -614
rect 928 -606 930 -596
rect 1243 -592 1263 -590
rect 1147 -606 1167 -604
rect 1147 -614 1167 -612
rect 791 -629 793 -619
rect 200 -661 220 -659
rect 200 -669 220 -667
rect 411 -671 441 -669
rect 411 -679 441 -677
rect 555 -669 580 -667
rect 555 -677 580 -675
rect 411 -687 441 -685
rect 109 -695 129 -693
rect 296 -695 316 -693
rect 109 -703 129 -701
rect 411 -695 441 -693
rect 296 -703 316 -701
rect 555 -685 580 -683
rect 683 -677 723 -675
rect 994 -673 1004 -671
rect 994 -681 1004 -679
rect 683 -685 723 -683
rect 555 -693 580 -691
rect 411 -703 441 -701
rect 473 -709 475 -699
rect 555 -701 580 -699
rect 606 -700 608 -690
rect 683 -693 723 -691
rect 994 -689 1004 -687
rect 994 -697 1004 -695
rect 683 -701 723 -699
rect 748 -709 750 -699
rect 994 -705 1004 -703
rect 411 -711 441 -709
rect 200 -717 220 -715
rect 1037 -711 1039 -701
rect 994 -713 1004 -711
rect 200 -725 220 -723
rect 91 -775 111 -773
rect 91 -783 111 -781
rect 136 -793 138 -783
<< ptransistor >>
rect 414 226 434 228
rect 414 218 434 220
rect 323 192 343 194
rect 510 192 530 194
rect 323 184 343 186
rect 510 184 530 186
rect 414 170 434 172
rect 414 162 434 164
rect 163 138 183 140
rect 163 130 183 132
rect 72 104 92 106
rect 259 104 279 106
rect 72 96 92 98
rect 259 96 279 98
rect 444 93 446 113
rect 572 93 574 113
rect 366 85 386 87
rect 163 82 183 84
rect 366 77 386 79
rect 484 84 524 86
rect 163 74 183 76
rect 484 76 524 78
rect 135 32 137 52
rect 57 24 77 26
rect 57 16 77 18
rect 367 7 369 27
rect 289 -1 309 1
rect 289 -9 309 -7
rect 413 2 473 4
rect 520 0 522 20
rect 413 -6 473 -4
rect 413 -14 473 -12
rect 162 -42 182 -40
rect 162 -50 182 -48
rect 71 -76 91 -74
rect 258 -76 278 -74
rect 71 -84 91 -82
rect 258 -84 278 -82
rect 372 -83 392 -81
rect 459 -86 461 -66
rect 372 -91 392 -89
rect 162 -98 182 -96
rect 372 -99 392 -97
rect 162 -106 182 -104
rect 134 -148 136 -128
rect 653 -129 673 -127
rect 653 -137 673 -135
rect 56 -156 76 -154
rect 56 -164 76 -162
rect 562 -163 582 -161
rect 294 -169 314 -167
rect 749 -163 769 -161
rect 562 -171 582 -169
rect 294 -177 314 -175
rect 749 -171 769 -169
rect 653 -185 673 -183
rect 653 -193 673 -191
rect 203 -203 223 -201
rect 390 -203 410 -201
rect 203 -211 223 -209
rect 390 -211 410 -209
rect 294 -225 314 -223
rect 294 -233 314 -231
rect 624 -259 626 -239
rect 546 -267 566 -265
rect 546 -275 566 -273
rect 162 -296 182 -294
rect 162 -304 182 -302
rect 377 -318 397 -316
rect 71 -330 91 -328
rect 474 -324 476 -304
rect 546 -320 566 -318
rect 377 -326 397 -324
rect 258 -330 278 -328
rect 71 -338 91 -336
rect 377 -334 397 -332
rect 258 -338 278 -336
rect 633 -323 635 -303
rect 693 -304 773 -302
rect 693 -312 773 -310
rect 821 -312 823 -292
rect 693 -320 773 -318
rect 546 -328 566 -326
rect 546 -336 566 -334
rect 377 -342 397 -340
rect 693 -328 773 -326
rect 162 -352 182 -350
rect 162 -360 182 -358
rect 801 -380 803 -360
rect 134 -402 136 -382
rect 723 -388 743 -386
rect 723 -396 743 -394
rect 56 -410 76 -408
rect 56 -418 76 -416
rect 305 -431 325 -429
rect 388 -436 390 -416
rect 441 -429 461 -427
rect 305 -439 325 -437
rect 305 -447 325 -445
rect 538 -435 540 -415
rect 587 -432 607 -430
rect 441 -437 461 -435
rect 441 -445 461 -443
rect 305 -455 325 -453
rect 305 -463 325 -461
rect 674 -435 676 -415
rect 587 -440 607 -438
rect 587 -448 607 -446
rect 441 -453 461 -451
rect 733 -452 833 -450
rect 879 -456 881 -436
rect 733 -460 833 -458
rect 733 -468 833 -466
rect 163 -478 183 -476
rect 733 -476 833 -474
rect 163 -486 183 -484
rect 733 -484 833 -482
rect 72 -512 92 -510
rect 259 -512 279 -510
rect 72 -520 92 -518
rect 259 -520 279 -518
rect 163 -534 183 -532
rect 163 -542 183 -540
rect 486 -547 506 -545
rect 1111 -550 1131 -548
rect 486 -555 506 -553
rect 1111 -558 1131 -556
rect 135 -584 137 -564
rect 395 -581 415 -579
rect 57 -592 77 -590
rect 57 -600 77 -598
rect 582 -581 602 -579
rect 928 -580 930 -560
rect 395 -589 415 -587
rect 582 -589 602 -587
rect 704 -600 724 -598
rect 486 -603 506 -601
rect 791 -603 793 -583
rect 850 -588 870 -586
rect 850 -596 870 -594
rect 1020 -584 1040 -582
rect 1207 -584 1227 -582
rect 1020 -592 1040 -590
rect 704 -608 724 -606
rect 486 -611 506 -609
rect 704 -616 724 -614
rect 1207 -592 1227 -590
rect 1111 -606 1131 -604
rect 1111 -614 1131 -612
rect 164 -661 184 -659
rect 164 -669 184 -667
rect 387 -671 397 -669
rect 387 -679 397 -677
rect 473 -683 475 -663
rect 523 -669 543 -667
rect 606 -674 608 -654
rect 523 -677 543 -675
rect 387 -687 397 -685
rect 73 -695 93 -693
rect 260 -695 280 -693
rect 73 -703 93 -701
rect 387 -695 397 -693
rect 260 -703 280 -701
rect 523 -685 543 -683
rect 651 -677 671 -675
rect 748 -683 750 -663
rect 862 -673 982 -671
rect 862 -681 982 -679
rect 651 -685 671 -683
rect 523 -693 543 -691
rect 387 -703 397 -701
rect 523 -701 543 -699
rect 651 -693 671 -691
rect 1037 -685 1039 -665
rect 862 -689 982 -687
rect 862 -697 982 -695
rect 651 -701 671 -699
rect 862 -705 982 -703
rect 387 -711 397 -709
rect 164 -717 184 -715
rect 862 -713 982 -711
rect 164 -725 184 -723
rect 136 -767 138 -747
rect 58 -775 78 -773
rect 58 -783 78 -781
<< ndiffusion >>
rect 450 228 470 229
rect 450 225 470 226
rect 450 220 470 221
rect 450 217 470 218
rect 359 194 379 195
rect 359 191 379 192
rect 546 194 566 195
rect 359 186 379 187
rect 359 183 379 184
rect 546 191 566 192
rect 546 186 566 187
rect 546 183 566 184
rect 450 172 470 173
rect 450 169 470 170
rect 450 164 470 165
rect 450 161 470 162
rect 199 140 219 141
rect 199 137 219 138
rect 199 132 219 133
rect 199 129 219 130
rect 108 106 128 107
rect 108 103 128 104
rect 295 106 315 107
rect 108 98 128 99
rect 108 95 128 96
rect 295 103 315 104
rect 295 98 315 99
rect 295 95 315 96
rect 199 84 219 85
rect 399 87 419 88
rect 199 81 219 82
rect 199 76 219 77
rect 399 84 419 85
rect 399 79 419 80
rect 536 86 546 87
rect 199 73 219 74
rect 399 76 419 77
rect 443 67 444 77
rect 446 67 447 77
rect 536 83 546 84
rect 536 78 546 79
rect 536 75 546 76
rect 571 67 572 77
rect 574 67 575 77
rect 90 26 110 27
rect 90 23 110 24
rect 90 18 110 19
rect 90 15 110 16
rect 134 6 135 16
rect 137 6 138 16
rect 322 1 342 2
rect 322 -2 342 -1
rect 322 -7 342 -6
rect 485 4 495 5
rect 485 1 495 2
rect 485 -4 495 -3
rect 322 -10 342 -9
rect 366 -19 367 -9
rect 369 -19 370 -9
rect 485 -7 495 -6
rect 485 -12 495 -11
rect 485 -15 495 -14
rect 519 -26 520 -16
rect 522 -26 523 -16
rect 198 -40 218 -39
rect 198 -43 218 -42
rect 198 -48 218 -47
rect 198 -51 218 -50
rect 107 -74 127 -73
rect 107 -77 127 -76
rect 294 -74 314 -73
rect 107 -82 127 -81
rect 107 -85 127 -84
rect 294 -77 314 -76
rect 294 -82 314 -81
rect 404 -81 434 -80
rect 294 -85 314 -84
rect 404 -84 434 -83
rect 404 -89 434 -88
rect 198 -96 218 -95
rect 198 -99 218 -98
rect 404 -92 434 -91
rect 404 -97 434 -96
rect 198 -104 218 -103
rect 404 -100 434 -99
rect 198 -107 218 -106
rect 458 -112 459 -102
rect 461 -112 462 -102
rect 689 -127 709 -126
rect 689 -130 709 -129
rect 689 -135 709 -134
rect 689 -138 709 -137
rect 89 -154 109 -153
rect 89 -157 109 -156
rect 89 -162 109 -161
rect 89 -165 109 -164
rect 133 -174 134 -164
rect 136 -174 137 -164
rect 598 -161 618 -160
rect 330 -167 350 -166
rect 330 -170 350 -169
rect 598 -164 618 -163
rect 785 -161 805 -160
rect 598 -169 618 -168
rect 330 -175 350 -174
rect 598 -172 618 -171
rect 785 -164 805 -163
rect 785 -169 805 -168
rect 785 -172 805 -171
rect 330 -178 350 -177
rect 689 -183 709 -182
rect 689 -186 709 -185
rect 689 -191 709 -190
rect 239 -201 259 -200
rect 239 -204 259 -203
rect 689 -194 709 -193
rect 426 -201 446 -200
rect 239 -209 259 -208
rect 239 -212 259 -211
rect 426 -204 446 -203
rect 426 -209 446 -208
rect 426 -212 446 -211
rect 330 -223 350 -222
rect 330 -226 350 -225
rect 330 -231 350 -230
rect 330 -234 350 -233
rect 579 -265 599 -264
rect 579 -268 599 -267
rect 579 -273 599 -272
rect 579 -276 599 -275
rect 623 -285 624 -275
rect 626 -285 627 -275
rect 198 -294 218 -293
rect 198 -297 218 -296
rect 198 -302 218 -301
rect 198 -305 218 -304
rect 409 -316 449 -315
rect 107 -328 127 -327
rect 107 -331 127 -330
rect 409 -319 449 -318
rect 409 -324 449 -323
rect 578 -318 608 -317
rect 294 -328 314 -327
rect 107 -336 127 -335
rect 107 -339 127 -338
rect 294 -331 314 -330
rect 409 -327 449 -326
rect 409 -332 449 -331
rect 294 -336 314 -335
rect 294 -339 314 -338
rect 409 -335 449 -334
rect 409 -340 449 -339
rect 578 -321 608 -320
rect 785 -302 795 -301
rect 785 -305 795 -304
rect 785 -310 795 -309
rect 785 -313 795 -312
rect 785 -318 795 -317
rect 578 -326 608 -325
rect 578 -329 608 -328
rect 578 -334 608 -333
rect 409 -343 449 -342
rect 198 -350 218 -349
rect 473 -350 474 -340
rect 476 -350 477 -340
rect 578 -337 608 -336
rect 785 -321 795 -320
rect 785 -326 795 -325
rect 785 -329 795 -328
rect 820 -338 821 -328
rect 823 -338 824 -328
rect 632 -349 633 -339
rect 635 -349 636 -339
rect 198 -353 218 -352
rect 198 -358 218 -357
rect 198 -361 218 -360
rect 756 -386 776 -385
rect 756 -389 776 -388
rect 756 -394 776 -393
rect 756 -397 776 -396
rect 89 -408 109 -407
rect 89 -411 109 -410
rect 89 -416 109 -415
rect 800 -406 801 -396
rect 803 -406 804 -396
rect 89 -419 109 -418
rect 133 -428 134 -418
rect 136 -428 137 -418
rect 337 -429 362 -428
rect 337 -432 362 -431
rect 473 -427 513 -426
rect 337 -437 362 -436
rect 337 -440 362 -439
rect 337 -445 362 -444
rect 337 -448 362 -447
rect 473 -430 513 -429
rect 473 -435 513 -434
rect 619 -430 649 -429
rect 473 -438 513 -437
rect 473 -443 513 -442
rect 337 -453 362 -452
rect 337 -456 362 -455
rect 337 -461 362 -460
rect 387 -462 388 -452
rect 390 -462 391 -452
rect 473 -446 513 -445
rect 473 -451 513 -450
rect 619 -433 649 -432
rect 619 -438 649 -437
rect 619 -441 649 -440
rect 619 -446 649 -445
rect 473 -454 513 -453
rect 537 -461 538 -451
rect 540 -461 541 -451
rect 619 -449 649 -448
rect 673 -461 674 -451
rect 676 -461 677 -451
rect 845 -450 855 -449
rect 845 -453 855 -452
rect 845 -458 855 -457
rect 337 -464 362 -463
rect 845 -461 855 -460
rect 845 -466 855 -465
rect 199 -476 219 -475
rect 845 -469 855 -468
rect 845 -474 855 -473
rect 199 -479 219 -478
rect 199 -484 219 -483
rect 845 -477 855 -476
rect 845 -482 855 -481
rect 878 -482 879 -472
rect 881 -482 882 -472
rect 199 -487 219 -486
rect 845 -485 855 -484
rect 108 -510 128 -509
rect 108 -513 128 -512
rect 295 -510 315 -509
rect 108 -518 128 -517
rect 108 -521 128 -520
rect 295 -513 315 -512
rect 295 -518 315 -517
rect 295 -521 315 -520
rect 199 -532 219 -531
rect 199 -535 219 -534
rect 199 -540 219 -539
rect 199 -543 219 -542
rect 522 -545 542 -544
rect 522 -548 542 -547
rect 1147 -548 1167 -547
rect 522 -553 542 -552
rect 522 -556 542 -555
rect 1147 -551 1167 -550
rect 1147 -556 1167 -555
rect 431 -579 451 -578
rect 90 -590 110 -589
rect 90 -593 110 -592
rect 90 -598 110 -597
rect 431 -582 451 -581
rect 618 -579 638 -578
rect 1147 -559 1167 -558
rect 431 -587 451 -586
rect 431 -590 451 -589
rect 618 -582 638 -581
rect 618 -587 638 -586
rect 618 -590 638 -589
rect 90 -601 110 -600
rect 134 -610 135 -600
rect 137 -610 138 -600
rect 522 -601 542 -600
rect 736 -598 766 -597
rect 522 -604 542 -603
rect 522 -609 542 -608
rect 736 -601 766 -600
rect 883 -586 903 -585
rect 883 -589 903 -588
rect 883 -594 903 -593
rect 1056 -582 1076 -581
rect 1056 -585 1076 -584
rect 1243 -582 1263 -581
rect 1056 -590 1076 -589
rect 883 -597 903 -596
rect 736 -606 766 -605
rect 522 -612 542 -611
rect 736 -609 766 -608
rect 736 -614 766 -613
rect 736 -617 766 -616
rect 927 -606 928 -596
rect 930 -606 931 -596
rect 1056 -593 1076 -592
rect 1243 -585 1263 -584
rect 1243 -590 1263 -589
rect 1243 -593 1263 -592
rect 1147 -604 1167 -603
rect 1147 -607 1167 -606
rect 1147 -612 1167 -611
rect 1147 -615 1167 -614
rect 790 -629 791 -619
rect 793 -629 794 -619
rect 200 -659 220 -658
rect 200 -662 220 -661
rect 200 -667 220 -666
rect 200 -670 220 -669
rect 411 -669 441 -668
rect 411 -672 441 -671
rect 411 -677 441 -676
rect 411 -680 441 -679
rect 555 -667 580 -666
rect 555 -670 580 -669
rect 555 -675 580 -674
rect 411 -685 441 -684
rect 109 -693 129 -692
rect 109 -696 129 -695
rect 296 -693 316 -692
rect 109 -701 129 -700
rect 109 -704 129 -703
rect 296 -696 316 -695
rect 411 -688 441 -687
rect 411 -693 441 -692
rect 296 -701 316 -700
rect 296 -704 316 -703
rect 411 -696 441 -695
rect 555 -678 580 -677
rect 555 -683 580 -682
rect 555 -686 580 -685
rect 683 -675 723 -674
rect 683 -678 723 -677
rect 683 -683 723 -682
rect 994 -671 1004 -670
rect 994 -674 1004 -673
rect 994 -679 1004 -678
rect 555 -691 580 -690
rect 411 -701 441 -700
rect 411 -704 441 -703
rect 411 -709 441 -708
rect 472 -709 473 -699
rect 475 -709 476 -699
rect 555 -694 580 -693
rect 555 -699 580 -698
rect 605 -700 606 -690
rect 608 -700 609 -690
rect 683 -686 723 -685
rect 683 -691 723 -690
rect 555 -702 580 -701
rect 683 -694 723 -693
rect 683 -699 723 -698
rect 994 -682 1004 -681
rect 994 -687 1004 -686
rect 994 -690 1004 -689
rect 994 -695 1004 -694
rect 683 -702 723 -701
rect 747 -709 748 -699
rect 750 -709 751 -699
rect 994 -698 1004 -697
rect 994 -703 1004 -702
rect 200 -715 220 -714
rect 411 -712 441 -711
rect 994 -706 1004 -705
rect 994 -711 1004 -710
rect 1036 -711 1037 -701
rect 1039 -711 1040 -701
rect 200 -718 220 -717
rect 994 -714 1004 -713
rect 200 -723 220 -722
rect 200 -726 220 -725
rect 91 -773 111 -772
rect 91 -776 111 -775
rect 91 -781 111 -780
rect 91 -784 111 -783
rect 135 -793 136 -783
rect 138 -793 139 -783
<< pdiffusion >>
rect 414 228 434 229
rect 414 225 434 226
rect 414 220 434 221
rect 414 217 434 218
rect 323 194 343 195
rect 323 191 343 192
rect 323 186 343 187
rect 510 194 530 195
rect 510 191 530 192
rect 323 183 343 184
rect 510 186 530 187
rect 510 183 530 184
rect 414 172 434 173
rect 414 169 434 170
rect 414 164 434 165
rect 414 161 434 162
rect 163 140 183 141
rect 163 137 183 138
rect 163 132 183 133
rect 163 129 183 130
rect 72 106 92 107
rect 72 103 92 104
rect 72 98 92 99
rect 259 106 279 107
rect 259 103 279 104
rect 72 95 92 96
rect 259 98 279 99
rect 259 95 279 96
rect 443 93 444 113
rect 446 93 447 113
rect 571 93 572 113
rect 574 93 575 113
rect 163 84 183 85
rect 366 87 386 88
rect 366 84 386 85
rect 163 81 183 82
rect 163 76 183 77
rect 366 79 386 80
rect 484 86 524 87
rect 484 83 524 84
rect 366 76 386 77
rect 163 73 183 74
rect 484 78 524 79
rect 484 75 524 76
rect 134 32 135 52
rect 137 32 138 52
rect 57 26 77 27
rect 57 23 77 24
rect 57 18 77 19
rect 57 15 77 16
rect 366 7 367 27
rect 369 7 370 27
rect 289 1 309 2
rect 289 -2 309 -1
rect 289 -7 309 -6
rect 413 4 473 5
rect 413 1 473 2
rect 413 -4 473 -3
rect 519 0 520 20
rect 522 0 523 20
rect 413 -7 473 -6
rect 289 -10 309 -9
rect 413 -12 473 -11
rect 413 -15 473 -14
rect 162 -40 182 -39
rect 162 -43 182 -42
rect 162 -48 182 -47
rect 162 -51 182 -50
rect 71 -74 91 -73
rect 71 -77 91 -76
rect 71 -82 91 -81
rect 258 -74 278 -73
rect 258 -77 278 -76
rect 71 -85 91 -84
rect 258 -82 278 -81
rect 372 -81 392 -80
rect 372 -84 392 -83
rect 258 -85 278 -84
rect 162 -96 182 -95
rect 372 -89 392 -88
rect 458 -86 459 -66
rect 461 -86 462 -66
rect 372 -92 392 -91
rect 162 -99 182 -98
rect 162 -104 182 -103
rect 372 -97 392 -96
rect 372 -100 392 -99
rect 162 -107 182 -106
rect 133 -148 134 -128
rect 136 -148 137 -128
rect 653 -127 673 -126
rect 653 -130 673 -129
rect 653 -135 673 -134
rect 653 -138 673 -137
rect 56 -154 76 -153
rect 56 -157 76 -156
rect 56 -162 76 -161
rect 56 -165 76 -164
rect 294 -167 314 -166
rect 562 -161 582 -160
rect 562 -164 582 -163
rect 294 -170 314 -169
rect 294 -175 314 -174
rect 562 -169 582 -168
rect 749 -161 769 -160
rect 749 -164 769 -163
rect 562 -172 582 -171
rect 749 -169 769 -168
rect 749 -172 769 -171
rect 294 -178 314 -177
rect 653 -183 673 -182
rect 653 -186 673 -185
rect 653 -191 673 -190
rect 653 -194 673 -193
rect 203 -201 223 -200
rect 203 -204 223 -203
rect 203 -209 223 -208
rect 390 -201 410 -200
rect 390 -204 410 -203
rect 203 -212 223 -211
rect 390 -209 410 -208
rect 390 -212 410 -211
rect 294 -223 314 -222
rect 294 -226 314 -225
rect 294 -231 314 -230
rect 294 -234 314 -233
rect 623 -259 624 -239
rect 626 -259 627 -239
rect 546 -265 566 -264
rect 546 -268 566 -267
rect 546 -273 566 -272
rect 546 -276 566 -275
rect 162 -294 182 -293
rect 162 -297 182 -296
rect 162 -302 182 -301
rect 162 -305 182 -304
rect 377 -316 397 -315
rect 377 -319 397 -318
rect 71 -328 91 -327
rect 71 -331 91 -330
rect 71 -336 91 -335
rect 258 -328 278 -327
rect 377 -324 397 -323
rect 473 -324 474 -304
rect 476 -324 477 -304
rect 546 -318 566 -317
rect 546 -321 566 -320
rect 377 -327 397 -326
rect 258 -331 278 -330
rect 71 -339 91 -338
rect 258 -336 278 -335
rect 377 -332 397 -331
rect 377 -335 397 -334
rect 258 -339 278 -338
rect 377 -340 397 -339
rect 546 -326 566 -325
rect 632 -323 633 -303
rect 635 -323 636 -303
rect 693 -302 773 -301
rect 693 -305 773 -304
rect 693 -310 773 -309
rect 820 -312 821 -292
rect 823 -312 824 -292
rect 693 -313 773 -312
rect 693 -318 773 -317
rect 693 -321 773 -320
rect 546 -329 566 -328
rect 546 -334 566 -333
rect 546 -337 566 -336
rect 377 -343 397 -342
rect 162 -350 182 -349
rect 693 -326 773 -325
rect 693 -329 773 -328
rect 162 -353 182 -352
rect 162 -358 182 -357
rect 162 -361 182 -360
rect 800 -380 801 -360
rect 803 -380 804 -360
rect 133 -402 134 -382
rect 136 -402 137 -382
rect 723 -386 743 -385
rect 723 -389 743 -388
rect 723 -394 743 -393
rect 723 -397 743 -396
rect 56 -408 76 -407
rect 56 -411 76 -410
rect 56 -416 76 -415
rect 56 -419 76 -418
rect 305 -429 325 -428
rect 305 -432 325 -431
rect 305 -437 325 -436
rect 387 -436 388 -416
rect 390 -436 391 -416
rect 441 -427 461 -426
rect 441 -430 461 -429
rect 305 -440 325 -439
rect 305 -445 325 -444
rect 305 -448 325 -447
rect 305 -453 325 -452
rect 441 -435 461 -434
rect 537 -435 538 -415
rect 540 -435 541 -415
rect 587 -430 607 -429
rect 587 -433 607 -432
rect 441 -438 461 -437
rect 441 -443 461 -442
rect 441 -446 461 -445
rect 305 -456 325 -455
rect 305 -461 325 -460
rect 441 -451 461 -450
rect 587 -438 607 -437
rect 673 -435 674 -415
rect 676 -435 677 -415
rect 587 -441 607 -440
rect 587 -446 607 -445
rect 587 -449 607 -448
rect 441 -454 461 -453
rect 733 -450 833 -449
rect 733 -453 833 -452
rect 733 -458 833 -457
rect 878 -456 879 -436
rect 881 -456 882 -436
rect 733 -461 833 -460
rect 305 -464 325 -463
rect 733 -466 833 -465
rect 733 -469 833 -468
rect 163 -476 183 -475
rect 733 -474 833 -473
rect 733 -477 833 -476
rect 163 -479 183 -478
rect 163 -484 183 -483
rect 733 -482 833 -481
rect 733 -485 833 -484
rect 163 -487 183 -486
rect 72 -510 92 -509
rect 72 -513 92 -512
rect 72 -518 92 -517
rect 259 -510 279 -509
rect 259 -513 279 -512
rect 72 -521 92 -520
rect 259 -518 279 -517
rect 259 -521 279 -520
rect 163 -532 183 -531
rect 163 -535 183 -534
rect 163 -540 183 -539
rect 163 -543 183 -542
rect 486 -545 506 -544
rect 486 -548 506 -547
rect 486 -553 506 -552
rect 1111 -548 1131 -547
rect 1111 -551 1131 -550
rect 486 -556 506 -555
rect 1111 -556 1131 -555
rect 1111 -559 1131 -558
rect 134 -584 135 -564
rect 137 -584 138 -564
rect 395 -579 415 -578
rect 395 -582 415 -581
rect 57 -590 77 -589
rect 57 -593 77 -592
rect 57 -598 77 -597
rect 395 -587 415 -586
rect 582 -579 602 -578
rect 927 -580 928 -560
rect 930 -580 931 -560
rect 582 -582 602 -581
rect 395 -590 415 -589
rect 582 -587 602 -586
rect 582 -590 602 -589
rect 57 -601 77 -600
rect 486 -601 506 -600
rect 704 -598 724 -597
rect 704 -601 724 -600
rect 486 -604 506 -603
rect 486 -609 506 -608
rect 704 -606 724 -605
rect 790 -603 791 -583
rect 793 -603 794 -583
rect 850 -586 870 -585
rect 850 -589 870 -588
rect 850 -594 870 -593
rect 1020 -582 1040 -581
rect 1020 -585 1040 -584
rect 1020 -590 1040 -589
rect 1207 -582 1227 -581
rect 1207 -585 1227 -584
rect 1020 -593 1040 -592
rect 850 -597 870 -596
rect 704 -609 724 -608
rect 486 -612 506 -611
rect 704 -614 724 -613
rect 704 -617 724 -616
rect 1207 -590 1227 -589
rect 1207 -593 1227 -592
rect 1111 -604 1131 -603
rect 1111 -607 1131 -606
rect 1111 -612 1131 -611
rect 1111 -615 1131 -614
rect 164 -659 184 -658
rect 164 -662 184 -661
rect 164 -667 184 -666
rect 164 -670 184 -669
rect 387 -669 397 -668
rect 387 -672 397 -671
rect 387 -677 397 -676
rect 387 -680 397 -679
rect 387 -685 397 -684
rect 472 -683 473 -663
rect 475 -683 476 -663
rect 523 -667 543 -666
rect 523 -670 543 -669
rect 523 -675 543 -674
rect 605 -674 606 -654
rect 608 -674 609 -654
rect 523 -678 543 -677
rect 387 -688 397 -687
rect 73 -693 93 -692
rect 73 -696 93 -695
rect 73 -701 93 -700
rect 260 -693 280 -692
rect 260 -696 280 -695
rect 73 -704 93 -703
rect 260 -701 280 -700
rect 387 -693 397 -692
rect 387 -696 397 -695
rect 260 -704 280 -703
rect 387 -701 397 -700
rect 523 -683 543 -682
rect 523 -686 543 -685
rect 523 -691 543 -690
rect 651 -675 671 -674
rect 651 -678 671 -677
rect 651 -683 671 -682
rect 747 -683 748 -663
rect 750 -683 751 -663
rect 862 -671 982 -670
rect 862 -674 982 -673
rect 862 -679 982 -678
rect 862 -682 982 -681
rect 651 -686 671 -685
rect 523 -694 543 -693
rect 387 -704 397 -703
rect 164 -715 184 -714
rect 387 -709 397 -708
rect 523 -699 543 -698
rect 651 -691 671 -690
rect 651 -694 671 -693
rect 523 -702 543 -701
rect 651 -699 671 -698
rect 862 -687 982 -686
rect 1036 -685 1037 -665
rect 1039 -685 1040 -665
rect 862 -690 982 -689
rect 862 -695 982 -694
rect 862 -698 982 -697
rect 651 -702 671 -701
rect 862 -703 982 -702
rect 862 -706 982 -705
rect 387 -712 397 -711
rect 862 -711 982 -710
rect 862 -714 982 -713
rect 164 -718 184 -717
rect 164 -723 184 -722
rect 164 -726 184 -725
rect 135 -767 136 -747
rect 138 -767 139 -747
rect 58 -773 78 -772
rect 58 -776 78 -775
rect 58 -781 78 -780
rect 58 -784 78 -783
<< ndcontact >>
rect 450 229 470 233
rect 450 221 470 225
rect 450 213 470 217
rect 359 195 379 199
rect 546 195 566 199
rect 359 187 379 191
rect 546 187 566 191
rect 359 179 379 183
rect 546 179 566 183
rect 450 173 470 177
rect 450 165 470 169
rect 450 157 470 161
rect 199 141 219 145
rect 199 133 219 137
rect 199 125 219 129
rect 108 107 128 111
rect 295 107 315 111
rect 108 99 128 103
rect 295 99 315 103
rect 108 91 128 95
rect 295 91 315 95
rect 199 85 219 89
rect 399 88 419 92
rect 199 77 219 81
rect 399 80 419 84
rect 536 87 546 91
rect 199 69 219 73
rect 399 72 419 76
rect 439 67 443 77
rect 447 67 451 77
rect 536 79 546 83
rect 536 71 546 75
rect 567 67 571 77
rect 575 67 579 77
rect 90 27 110 31
rect 90 19 110 23
rect 90 11 110 15
rect 130 6 134 16
rect 138 6 142 16
rect 322 2 342 6
rect 322 -6 342 -2
rect 485 5 495 9
rect 485 -3 495 1
rect 322 -14 342 -10
rect 362 -19 366 -9
rect 370 -19 374 -9
rect 485 -11 495 -7
rect 485 -19 495 -15
rect 515 -26 519 -16
rect 523 -26 527 -16
rect 198 -39 218 -35
rect 198 -47 218 -43
rect 198 -55 218 -51
rect 107 -73 127 -69
rect 294 -73 314 -69
rect 107 -81 127 -77
rect 294 -81 314 -77
rect 404 -80 434 -76
rect 107 -89 127 -85
rect 294 -89 314 -85
rect 198 -95 218 -91
rect 404 -88 434 -84
rect 198 -103 218 -99
rect 404 -96 434 -92
rect 404 -104 434 -100
rect 198 -111 218 -107
rect 454 -112 458 -102
rect 462 -112 466 -102
rect 689 -126 709 -122
rect 689 -134 709 -130
rect 689 -142 709 -138
rect 89 -153 109 -149
rect 89 -161 109 -157
rect 89 -169 109 -165
rect 129 -174 133 -164
rect 137 -174 141 -164
rect 330 -166 350 -162
rect 598 -160 618 -156
rect 330 -174 350 -170
rect 785 -160 805 -156
rect 598 -168 618 -164
rect 785 -168 805 -164
rect 598 -176 618 -172
rect 785 -176 805 -172
rect 330 -182 350 -178
rect 689 -182 709 -178
rect 689 -190 709 -186
rect 239 -200 259 -196
rect 426 -200 446 -196
rect 689 -198 709 -194
rect 239 -208 259 -204
rect 426 -208 446 -204
rect 239 -216 259 -212
rect 426 -216 446 -212
rect 330 -222 350 -218
rect 330 -230 350 -226
rect 330 -238 350 -234
rect 579 -264 599 -260
rect 579 -272 599 -268
rect 579 -280 599 -276
rect 619 -285 623 -275
rect 627 -285 631 -275
rect 198 -293 218 -289
rect 198 -301 218 -297
rect 198 -309 218 -305
rect 409 -315 449 -311
rect 107 -327 127 -323
rect 294 -327 314 -323
rect 409 -323 449 -319
rect 578 -317 608 -313
rect 107 -335 127 -331
rect 294 -335 314 -331
rect 409 -331 449 -327
rect 107 -343 127 -339
rect 294 -343 314 -339
rect 409 -339 449 -335
rect 578 -325 608 -321
rect 785 -301 795 -297
rect 785 -309 795 -305
rect 785 -317 795 -313
rect 578 -333 608 -329
rect 198 -349 218 -345
rect 409 -347 449 -343
rect 469 -350 473 -340
rect 477 -350 481 -340
rect 578 -341 608 -337
rect 785 -325 795 -321
rect 785 -333 795 -329
rect 816 -338 820 -328
rect 824 -338 828 -328
rect 628 -349 632 -339
rect 636 -349 640 -339
rect 198 -357 218 -353
rect 198 -365 218 -361
rect 756 -385 776 -381
rect 756 -393 776 -389
rect 756 -401 776 -397
rect 89 -407 109 -403
rect 89 -415 109 -411
rect 796 -406 800 -396
rect 804 -406 808 -396
rect 89 -423 109 -419
rect 129 -428 133 -418
rect 137 -428 141 -418
rect 337 -428 362 -424
rect 337 -436 362 -432
rect 473 -426 513 -422
rect 337 -444 362 -440
rect 337 -452 362 -448
rect 473 -434 513 -430
rect 619 -429 649 -425
rect 473 -442 513 -438
rect 337 -460 362 -456
rect 383 -462 387 -452
rect 391 -462 395 -452
rect 473 -450 513 -446
rect 619 -437 649 -433
rect 619 -445 649 -441
rect 473 -458 513 -454
rect 533 -461 537 -451
rect 541 -461 545 -451
rect 619 -453 649 -449
rect 669 -461 673 -451
rect 677 -461 681 -451
rect 845 -449 855 -445
rect 845 -457 855 -453
rect 337 -468 362 -464
rect 845 -465 855 -461
rect 199 -475 219 -471
rect 845 -473 855 -469
rect 199 -483 219 -479
rect 845 -481 855 -477
rect 874 -482 878 -472
rect 882 -482 886 -472
rect 199 -491 219 -487
rect 845 -489 855 -485
rect 108 -509 128 -505
rect 295 -509 315 -505
rect 108 -517 128 -513
rect 295 -517 315 -513
rect 108 -525 128 -521
rect 295 -525 315 -521
rect 199 -531 219 -527
rect 199 -539 219 -535
rect 199 -547 219 -543
rect 522 -544 542 -540
rect 522 -552 542 -548
rect 1147 -547 1167 -543
rect 522 -560 542 -556
rect 1147 -555 1167 -551
rect 431 -578 451 -574
rect 90 -589 110 -585
rect 90 -597 110 -593
rect 618 -578 638 -574
rect 1147 -563 1167 -559
rect 431 -586 451 -582
rect 618 -586 638 -582
rect 431 -594 451 -590
rect 618 -594 638 -590
rect 90 -605 110 -601
rect 130 -610 134 -600
rect 138 -610 142 -600
rect 522 -600 542 -596
rect 736 -597 766 -593
rect 522 -608 542 -604
rect 736 -605 766 -601
rect 883 -585 903 -581
rect 883 -593 903 -589
rect 1056 -581 1076 -577
rect 1243 -581 1263 -577
rect 1056 -589 1076 -585
rect 883 -601 903 -597
rect 522 -616 542 -612
rect 736 -613 766 -609
rect 736 -621 766 -617
rect 923 -606 927 -596
rect 931 -606 935 -596
rect 1243 -589 1263 -585
rect 1056 -597 1076 -593
rect 1243 -597 1263 -593
rect 1147 -603 1167 -599
rect 1147 -611 1167 -607
rect 1147 -619 1167 -615
rect 786 -629 790 -619
rect 794 -629 798 -619
rect 200 -658 220 -654
rect 200 -666 220 -662
rect 200 -674 220 -670
rect 411 -668 441 -664
rect 411 -676 441 -672
rect 411 -684 441 -680
rect 555 -666 580 -662
rect 555 -674 580 -670
rect 109 -692 129 -688
rect 296 -692 316 -688
rect 109 -700 129 -696
rect 411 -692 441 -688
rect 296 -700 316 -696
rect 109 -708 129 -704
rect 411 -700 441 -696
rect 555 -682 580 -678
rect 555 -690 580 -686
rect 683 -674 723 -670
rect 683 -682 723 -678
rect 994 -670 1004 -666
rect 994 -678 1004 -674
rect 296 -708 316 -704
rect 200 -714 220 -710
rect 411 -708 441 -704
rect 468 -709 472 -699
rect 476 -709 480 -699
rect 555 -698 580 -694
rect 601 -700 605 -690
rect 609 -700 613 -690
rect 683 -690 723 -686
rect 555 -706 580 -702
rect 683 -698 723 -694
rect 994 -686 1004 -682
rect 994 -694 1004 -690
rect 683 -706 723 -702
rect 743 -709 747 -699
rect 751 -709 755 -699
rect 994 -702 1004 -698
rect 411 -716 441 -712
rect 994 -710 1004 -706
rect 1032 -711 1036 -701
rect 1040 -711 1044 -701
rect 994 -718 1004 -714
rect 200 -722 220 -718
rect 200 -730 220 -726
rect 91 -772 111 -768
rect 91 -780 111 -776
rect 91 -788 111 -784
rect 131 -793 135 -783
rect 139 -793 143 -783
<< pdcontact >>
rect 414 229 434 233
rect 414 221 434 225
rect 414 213 434 217
rect 323 195 343 199
rect 510 195 530 199
rect 323 187 343 191
rect 510 187 530 191
rect 323 179 343 183
rect 510 179 530 183
rect 414 173 434 177
rect 414 165 434 169
rect 414 157 434 161
rect 163 141 183 145
rect 163 133 183 137
rect 163 125 183 129
rect 72 107 92 111
rect 259 107 279 111
rect 72 99 92 103
rect 259 99 279 103
rect 72 91 92 95
rect 259 91 279 95
rect 439 93 443 113
rect 447 93 451 113
rect 567 93 571 113
rect 575 93 579 113
rect 163 85 183 89
rect 366 88 386 92
rect 163 77 183 81
rect 366 80 386 84
rect 484 87 524 91
rect 484 79 524 83
rect 163 69 183 73
rect 366 72 386 76
rect 484 71 524 75
rect 130 32 134 52
rect 138 32 142 52
rect 57 27 77 31
rect 57 19 77 23
rect 57 11 77 15
rect 362 7 366 27
rect 370 7 374 27
rect 289 2 309 6
rect 289 -6 309 -2
rect 413 5 473 9
rect 413 -3 473 1
rect 515 0 519 20
rect 523 0 527 20
rect 289 -14 309 -10
rect 413 -11 473 -7
rect 413 -19 473 -15
rect 162 -39 182 -35
rect 162 -47 182 -43
rect 162 -55 182 -51
rect 71 -73 91 -69
rect 258 -73 278 -69
rect 71 -81 91 -77
rect 258 -81 278 -77
rect 71 -89 91 -85
rect 372 -80 392 -76
rect 258 -89 278 -85
rect 372 -88 392 -84
rect 162 -95 182 -91
rect 454 -86 458 -66
rect 462 -86 466 -66
rect 372 -96 392 -92
rect 162 -103 182 -99
rect 372 -104 392 -100
rect 162 -111 182 -107
rect 653 -126 673 -122
rect 129 -148 133 -128
rect 137 -148 141 -128
rect 653 -134 673 -130
rect 653 -142 673 -138
rect 56 -153 76 -149
rect 56 -161 76 -157
rect 562 -160 582 -156
rect 56 -169 76 -165
rect 294 -166 314 -162
rect 749 -160 769 -156
rect 562 -168 582 -164
rect 294 -174 314 -170
rect 749 -168 769 -164
rect 562 -176 582 -172
rect 749 -176 769 -172
rect 294 -182 314 -178
rect 653 -182 673 -178
rect 653 -190 673 -186
rect 203 -200 223 -196
rect 390 -200 410 -196
rect 203 -208 223 -204
rect 653 -198 673 -194
rect 390 -208 410 -204
rect 203 -216 223 -212
rect 390 -216 410 -212
rect 294 -222 314 -218
rect 294 -230 314 -226
rect 294 -238 314 -234
rect 619 -259 623 -239
rect 627 -259 631 -239
rect 546 -264 566 -260
rect 546 -272 566 -268
rect 546 -280 566 -276
rect 162 -293 182 -289
rect 162 -301 182 -297
rect 693 -301 773 -297
rect 162 -309 182 -305
rect 377 -315 397 -311
rect 377 -323 397 -319
rect 71 -327 91 -323
rect 258 -327 278 -323
rect 71 -335 91 -331
rect 469 -324 473 -304
rect 477 -324 481 -304
rect 546 -317 566 -313
rect 258 -335 278 -331
rect 71 -343 91 -339
rect 377 -331 397 -327
rect 258 -343 278 -339
rect 377 -339 397 -335
rect 546 -325 566 -321
rect 628 -323 632 -303
rect 636 -323 640 -303
rect 693 -309 773 -305
rect 816 -312 820 -292
rect 824 -312 828 -292
rect 693 -317 773 -313
rect 546 -333 566 -329
rect 162 -349 182 -345
rect 377 -347 397 -343
rect 546 -341 566 -337
rect 693 -325 773 -321
rect 693 -333 773 -329
rect 162 -357 182 -353
rect 162 -365 182 -361
rect 796 -380 800 -360
rect 804 -380 808 -360
rect 129 -402 133 -382
rect 137 -402 141 -382
rect 723 -385 743 -381
rect 723 -393 743 -389
rect 723 -401 743 -397
rect 56 -407 76 -403
rect 56 -415 76 -411
rect 56 -423 76 -419
rect 305 -428 325 -424
rect 305 -436 325 -432
rect 383 -436 387 -416
rect 391 -436 395 -416
rect 441 -426 461 -422
rect 441 -434 461 -430
rect 305 -444 325 -440
rect 305 -452 325 -448
rect 533 -435 537 -415
rect 541 -435 545 -415
rect 587 -429 607 -425
rect 441 -442 461 -438
rect 441 -450 461 -446
rect 305 -460 325 -456
rect 587 -437 607 -433
rect 669 -435 673 -415
rect 677 -435 681 -415
rect 587 -445 607 -441
rect 441 -458 461 -454
rect 587 -453 607 -449
rect 733 -449 833 -445
rect 733 -457 833 -453
rect 874 -456 878 -436
rect 882 -456 886 -436
rect 305 -468 325 -464
rect 733 -465 833 -461
rect 163 -475 183 -471
rect 733 -473 833 -469
rect 163 -483 183 -479
rect 733 -481 833 -477
rect 163 -491 183 -487
rect 733 -489 833 -485
rect 72 -509 92 -505
rect 259 -509 279 -505
rect 72 -517 92 -513
rect 259 -517 279 -513
rect 72 -525 92 -521
rect 259 -525 279 -521
rect 163 -531 183 -527
rect 163 -539 183 -535
rect 163 -547 183 -543
rect 486 -544 506 -540
rect 1111 -547 1131 -543
rect 486 -552 506 -548
rect 1111 -555 1131 -551
rect 486 -560 506 -556
rect 130 -584 134 -564
rect 138 -584 142 -564
rect 395 -578 415 -574
rect 582 -578 602 -574
rect 57 -589 77 -585
rect 57 -597 77 -593
rect 395 -586 415 -582
rect 923 -580 927 -560
rect 931 -580 935 -560
rect 1111 -563 1131 -559
rect 582 -586 602 -582
rect 395 -594 415 -590
rect 582 -594 602 -590
rect 486 -600 506 -596
rect 57 -605 77 -601
rect 704 -597 724 -593
rect 486 -608 506 -604
rect 704 -605 724 -601
rect 786 -603 790 -583
rect 794 -603 798 -583
rect 850 -585 870 -581
rect 850 -593 870 -589
rect 1020 -581 1040 -577
rect 1207 -581 1227 -577
rect 1020 -589 1040 -585
rect 1207 -589 1227 -585
rect 850 -601 870 -597
rect 486 -616 506 -612
rect 704 -613 724 -609
rect 704 -621 724 -617
rect 1020 -597 1040 -593
rect 1207 -597 1227 -593
rect 1111 -603 1131 -599
rect 1111 -611 1131 -607
rect 1111 -619 1131 -615
rect 164 -658 184 -654
rect 164 -666 184 -662
rect 387 -668 397 -664
rect 164 -674 184 -670
rect 387 -676 397 -672
rect 387 -684 397 -680
rect 468 -683 472 -663
rect 476 -683 480 -663
rect 523 -666 543 -662
rect 523 -674 543 -670
rect 601 -674 605 -654
rect 609 -674 613 -654
rect 651 -674 671 -670
rect 523 -682 543 -678
rect 73 -692 93 -688
rect 260 -692 280 -688
rect 73 -700 93 -696
rect 387 -692 397 -688
rect 260 -700 280 -696
rect 73 -708 93 -704
rect 387 -700 397 -696
rect 260 -708 280 -704
rect 523 -690 543 -686
rect 651 -682 671 -678
rect 743 -683 747 -663
rect 751 -683 755 -663
rect 862 -670 982 -666
rect 862 -678 982 -674
rect 651 -690 671 -686
rect 523 -698 543 -694
rect 387 -708 397 -704
rect 164 -714 184 -710
rect 651 -698 671 -694
rect 523 -706 543 -702
rect 862 -686 982 -682
rect 1032 -685 1036 -665
rect 1040 -685 1044 -665
rect 862 -694 982 -690
rect 651 -706 671 -702
rect 862 -702 982 -698
rect 387 -716 397 -712
rect 862 -710 982 -706
rect 164 -722 184 -718
rect 862 -718 982 -714
rect 164 -730 184 -726
rect 131 -767 135 -747
rect 139 -767 143 -747
rect 58 -772 78 -768
rect 58 -780 78 -776
rect 58 -788 78 -784
<< polysilicon >>
rect 402 226 414 228
rect 434 226 450 228
rect 470 226 473 228
rect 402 218 414 220
rect 434 218 450 220
rect 470 218 473 220
rect 311 192 323 194
rect 343 192 359 194
rect 379 192 382 194
rect 498 192 510 194
rect 530 192 546 194
rect 566 192 569 194
rect 311 184 323 186
rect 343 184 359 186
rect 379 184 382 186
rect 498 184 510 186
rect 530 184 546 186
rect 566 184 569 186
rect 402 170 414 172
rect 434 170 450 172
rect 470 170 473 172
rect 402 162 414 164
rect 434 162 450 164
rect 470 162 473 164
rect 151 138 163 140
rect 183 138 199 140
rect 219 138 222 140
rect 151 130 163 132
rect 183 130 199 132
rect 219 130 222 132
rect 444 113 446 116
rect 572 113 574 116
rect 60 104 72 106
rect 92 104 108 106
rect 128 104 131 106
rect 247 104 259 106
rect 279 104 295 106
rect 315 104 318 106
rect 60 96 72 98
rect 92 96 108 98
rect 128 96 131 98
rect 247 96 259 98
rect 279 96 295 98
rect 315 96 318 98
rect 357 85 366 87
rect 386 85 399 87
rect 419 85 422 87
rect 151 82 163 84
rect 183 82 199 84
rect 219 82 222 84
rect 357 77 366 79
rect 386 77 399 79
rect 419 77 422 79
rect 444 77 446 93
rect 475 84 484 86
rect 524 84 536 86
rect 546 84 549 86
rect 151 74 163 76
rect 183 74 199 76
rect 219 74 222 76
rect 475 76 484 78
rect 524 76 536 78
rect 546 76 549 78
rect 572 77 574 93
rect 444 64 446 67
rect 572 64 574 67
rect 135 52 137 55
rect 48 24 57 26
rect 77 24 90 26
rect 110 24 113 26
rect 48 16 57 18
rect 77 16 90 18
rect 110 16 113 18
rect 135 16 137 32
rect 367 27 369 30
rect 520 20 522 23
rect 135 3 137 6
rect 280 -1 289 1
rect 309 -1 322 1
rect 342 -1 345 1
rect 280 -9 289 -7
rect 309 -9 322 -7
rect 342 -9 345 -7
rect 367 -9 369 7
rect 404 2 413 4
rect 473 2 485 4
rect 495 2 498 4
rect 404 -6 413 -4
rect 473 -6 485 -4
rect 495 -6 498 -4
rect 404 -14 413 -12
rect 473 -14 485 -12
rect 495 -14 498 -12
rect 520 -16 522 0
rect 367 -22 369 -19
rect 520 -29 522 -26
rect 150 -42 162 -40
rect 182 -42 198 -40
rect 218 -42 221 -40
rect 150 -50 162 -48
rect 182 -50 198 -48
rect 218 -50 221 -48
rect 459 -66 461 -63
rect 59 -76 71 -74
rect 91 -76 107 -74
rect 127 -76 130 -74
rect 246 -76 258 -74
rect 278 -76 294 -74
rect 314 -76 317 -74
rect 59 -84 71 -82
rect 91 -84 107 -82
rect 127 -84 130 -82
rect 246 -84 258 -82
rect 278 -84 294 -82
rect 314 -84 317 -82
rect 363 -83 372 -81
rect 392 -83 404 -81
rect 434 -83 437 -81
rect 363 -91 372 -89
rect 392 -91 404 -89
rect 434 -91 437 -89
rect 150 -98 162 -96
rect 182 -98 198 -96
rect 218 -98 221 -96
rect 363 -99 372 -97
rect 392 -99 404 -97
rect 434 -99 437 -97
rect 459 -102 461 -86
rect 150 -106 162 -104
rect 182 -106 198 -104
rect 218 -106 221 -104
rect 459 -115 461 -112
rect 134 -128 136 -125
rect 641 -129 653 -127
rect 673 -129 689 -127
rect 709 -129 712 -127
rect 641 -137 653 -135
rect 673 -137 689 -135
rect 709 -137 712 -135
rect 47 -156 56 -154
rect 76 -156 89 -154
rect 109 -156 112 -154
rect 47 -164 56 -162
rect 76 -164 89 -162
rect 109 -164 112 -162
rect 134 -164 136 -148
rect 550 -163 562 -161
rect 582 -163 598 -161
rect 618 -163 621 -161
rect 282 -169 294 -167
rect 314 -169 330 -167
rect 350 -169 353 -167
rect 134 -177 136 -174
rect 737 -163 749 -161
rect 769 -163 785 -161
rect 805 -163 808 -161
rect 550 -171 562 -169
rect 582 -171 598 -169
rect 618 -171 621 -169
rect 282 -177 294 -175
rect 314 -177 330 -175
rect 350 -177 353 -175
rect 737 -171 749 -169
rect 769 -171 785 -169
rect 805 -171 808 -169
rect 641 -185 653 -183
rect 673 -185 689 -183
rect 709 -185 712 -183
rect 641 -193 653 -191
rect 673 -193 689 -191
rect 709 -193 712 -191
rect 191 -203 203 -201
rect 223 -203 239 -201
rect 259 -203 262 -201
rect 378 -203 390 -201
rect 410 -203 426 -201
rect 446 -203 449 -201
rect 191 -211 203 -209
rect 223 -211 239 -209
rect 259 -211 262 -209
rect 378 -211 390 -209
rect 410 -211 426 -209
rect 446 -211 449 -209
rect 282 -225 294 -223
rect 314 -225 330 -223
rect 350 -225 353 -223
rect 282 -233 294 -231
rect 314 -233 330 -231
rect 350 -233 353 -231
rect 624 -239 626 -236
rect 537 -267 546 -265
rect 566 -267 579 -265
rect 599 -267 602 -265
rect 537 -275 546 -273
rect 566 -275 579 -273
rect 599 -275 602 -273
rect 624 -275 626 -259
rect 624 -288 626 -285
rect 821 -292 823 -289
rect 150 -296 162 -294
rect 182 -296 198 -294
rect 218 -296 221 -294
rect 150 -304 162 -302
rect 182 -304 198 -302
rect 218 -304 221 -302
rect 474 -304 476 -301
rect 633 -303 635 -300
rect 368 -318 377 -316
rect 397 -318 409 -316
rect 449 -318 452 -316
rect 59 -330 71 -328
rect 91 -330 107 -328
rect 127 -330 130 -328
rect 537 -320 546 -318
rect 566 -320 578 -318
rect 608 -320 611 -318
rect 368 -326 377 -324
rect 397 -326 409 -324
rect 449 -326 452 -324
rect 246 -330 258 -328
rect 278 -330 294 -328
rect 314 -330 317 -328
rect 59 -338 71 -336
rect 91 -338 107 -336
rect 127 -338 130 -336
rect 368 -334 377 -332
rect 397 -334 409 -332
rect 449 -334 452 -332
rect 246 -338 258 -336
rect 278 -338 294 -336
rect 314 -338 317 -336
rect 474 -340 476 -324
rect 684 -304 693 -302
rect 773 -304 785 -302
rect 795 -304 798 -302
rect 684 -312 693 -310
rect 773 -312 785 -310
rect 795 -312 798 -310
rect 684 -320 693 -318
rect 773 -320 785 -318
rect 795 -320 798 -318
rect 537 -328 546 -326
rect 566 -328 578 -326
rect 608 -328 611 -326
rect 537 -336 546 -334
rect 566 -336 578 -334
rect 608 -336 611 -334
rect 368 -342 377 -340
rect 397 -342 409 -340
rect 449 -342 452 -340
rect 633 -339 635 -323
rect 684 -328 693 -326
rect 773 -328 785 -326
rect 795 -328 798 -326
rect 821 -328 823 -312
rect 821 -341 823 -338
rect 150 -352 162 -350
rect 182 -352 198 -350
rect 218 -352 221 -350
rect 474 -353 476 -350
rect 633 -352 635 -349
rect 150 -360 162 -358
rect 182 -360 198 -358
rect 218 -360 221 -358
rect 801 -360 803 -357
rect 134 -382 136 -379
rect 714 -388 723 -386
rect 743 -388 756 -386
rect 776 -388 779 -386
rect 714 -396 723 -394
rect 743 -396 756 -394
rect 776 -396 779 -394
rect 801 -396 803 -380
rect 47 -410 56 -408
rect 76 -410 89 -408
rect 109 -410 112 -408
rect 47 -418 56 -416
rect 76 -418 89 -416
rect 109 -418 112 -416
rect 134 -418 136 -402
rect 801 -409 803 -406
rect 388 -416 390 -413
rect 538 -415 540 -412
rect 674 -415 676 -412
rect 134 -431 136 -428
rect 296 -431 305 -429
rect 325 -431 337 -429
rect 362 -431 365 -429
rect 432 -429 441 -427
rect 461 -429 473 -427
rect 513 -429 516 -427
rect 296 -439 305 -437
rect 325 -439 337 -437
rect 362 -439 365 -437
rect 296 -447 305 -445
rect 325 -447 337 -445
rect 362 -447 365 -445
rect 388 -452 390 -436
rect 578 -432 587 -430
rect 607 -432 619 -430
rect 649 -432 652 -430
rect 432 -437 441 -435
rect 461 -437 473 -435
rect 513 -437 516 -435
rect 432 -445 441 -443
rect 461 -445 473 -443
rect 513 -445 516 -443
rect 296 -455 305 -453
rect 325 -455 337 -453
rect 362 -455 375 -453
rect 373 -458 375 -455
rect 296 -463 305 -461
rect 325 -463 337 -461
rect 362 -463 365 -461
rect 538 -451 540 -435
rect 578 -440 587 -438
rect 607 -440 619 -438
rect 649 -440 652 -438
rect 578 -448 587 -446
rect 607 -448 619 -446
rect 649 -448 652 -446
rect 432 -453 441 -451
rect 461 -453 473 -451
rect 513 -453 516 -451
rect 674 -451 676 -435
rect 879 -436 881 -433
rect 724 -452 733 -450
rect 833 -452 845 -450
rect 855 -452 858 -450
rect 724 -460 733 -458
rect 833 -460 845 -458
rect 855 -460 858 -458
rect 388 -465 390 -462
rect 538 -464 540 -461
rect 674 -464 676 -461
rect 724 -468 733 -466
rect 833 -468 845 -466
rect 855 -468 858 -466
rect 151 -478 163 -476
rect 183 -478 199 -476
rect 219 -478 222 -476
rect 879 -472 881 -456
rect 724 -476 733 -474
rect 833 -476 845 -474
rect 855 -476 858 -474
rect 151 -486 163 -484
rect 183 -486 199 -484
rect 219 -486 222 -484
rect 724 -484 733 -482
rect 833 -484 845 -482
rect 855 -484 858 -482
rect 879 -485 881 -482
rect 60 -512 72 -510
rect 92 -512 108 -510
rect 128 -512 131 -510
rect 247 -512 259 -510
rect 279 -512 295 -510
rect 315 -512 318 -510
rect 60 -520 72 -518
rect 92 -520 108 -518
rect 128 -520 131 -518
rect 247 -520 259 -518
rect 279 -520 295 -518
rect 315 -520 318 -518
rect 151 -534 163 -532
rect 183 -534 199 -532
rect 219 -534 222 -532
rect 151 -542 163 -540
rect 183 -542 199 -540
rect 219 -542 222 -540
rect 474 -547 486 -545
rect 506 -547 522 -545
rect 542 -547 545 -545
rect 1099 -550 1111 -548
rect 1131 -550 1147 -548
rect 1167 -550 1170 -548
rect 474 -555 486 -553
rect 506 -555 522 -553
rect 542 -555 545 -553
rect 928 -560 930 -557
rect 1099 -558 1111 -556
rect 1131 -558 1147 -556
rect 1167 -558 1170 -556
rect 135 -564 137 -561
rect 383 -581 395 -579
rect 415 -581 431 -579
rect 451 -581 454 -579
rect 48 -592 57 -590
rect 77 -592 90 -590
rect 110 -592 113 -590
rect 48 -600 57 -598
rect 77 -600 90 -598
rect 110 -600 113 -598
rect 135 -600 137 -584
rect 570 -581 582 -579
rect 602 -581 618 -579
rect 638 -581 641 -579
rect 383 -589 395 -587
rect 415 -589 431 -587
rect 451 -589 454 -587
rect 791 -583 793 -580
rect 570 -589 582 -587
rect 602 -589 618 -587
rect 638 -589 641 -587
rect 695 -600 704 -598
rect 724 -600 736 -598
rect 766 -600 769 -598
rect 474 -603 486 -601
rect 506 -603 522 -601
rect 542 -603 545 -601
rect 135 -613 137 -610
rect 841 -588 850 -586
rect 870 -588 883 -586
rect 903 -588 906 -586
rect 841 -596 850 -594
rect 870 -596 883 -594
rect 903 -596 906 -594
rect 928 -596 930 -580
rect 1008 -584 1020 -582
rect 1040 -584 1056 -582
rect 1076 -584 1079 -582
rect 1195 -584 1207 -582
rect 1227 -584 1243 -582
rect 1263 -584 1266 -582
rect 1008 -592 1020 -590
rect 1040 -592 1056 -590
rect 1076 -592 1079 -590
rect 695 -608 704 -606
rect 724 -608 736 -606
rect 766 -608 769 -606
rect 474 -611 486 -609
rect 506 -611 522 -609
rect 542 -611 545 -609
rect 695 -616 704 -614
rect 724 -616 736 -614
rect 766 -616 769 -614
rect 791 -619 793 -603
rect 1195 -592 1207 -590
rect 1227 -592 1243 -590
rect 1263 -592 1266 -590
rect 928 -609 930 -606
rect 1099 -606 1111 -604
rect 1131 -606 1147 -604
rect 1167 -606 1170 -604
rect 1099 -614 1111 -612
rect 1131 -614 1147 -612
rect 1167 -614 1170 -612
rect 791 -632 793 -629
rect 606 -654 608 -651
rect 152 -661 164 -659
rect 184 -661 200 -659
rect 220 -661 223 -659
rect 473 -663 475 -660
rect 152 -669 164 -667
rect 184 -669 200 -667
rect 220 -669 223 -667
rect 377 -671 387 -669
rect 397 -671 411 -669
rect 441 -671 444 -669
rect 377 -679 387 -677
rect 397 -679 411 -677
rect 441 -679 444 -677
rect 514 -669 523 -667
rect 543 -669 555 -667
rect 580 -669 583 -667
rect 748 -663 750 -660
rect 514 -677 523 -675
rect 543 -677 555 -675
rect 580 -677 583 -675
rect 377 -687 387 -685
rect 397 -687 411 -685
rect 441 -687 444 -685
rect 61 -695 73 -693
rect 93 -695 109 -693
rect 129 -695 132 -693
rect 248 -695 260 -693
rect 280 -695 296 -693
rect 316 -695 319 -693
rect 61 -703 73 -701
rect 93 -703 109 -701
rect 129 -703 132 -701
rect 377 -695 387 -693
rect 397 -695 411 -693
rect 441 -695 444 -693
rect 248 -703 260 -701
rect 280 -703 296 -701
rect 316 -703 319 -701
rect 473 -699 475 -683
rect 514 -685 523 -683
rect 543 -685 555 -683
rect 580 -685 583 -683
rect 606 -690 608 -674
rect 642 -677 651 -675
rect 671 -677 683 -675
rect 723 -677 726 -675
rect 1037 -665 1039 -662
rect 851 -673 862 -671
rect 982 -673 994 -671
rect 1004 -673 1007 -671
rect 851 -681 862 -679
rect 982 -681 994 -679
rect 1004 -681 1007 -679
rect 642 -685 651 -683
rect 671 -685 683 -683
rect 723 -685 726 -683
rect 514 -693 523 -691
rect 543 -693 555 -691
rect 580 -693 595 -691
rect 377 -703 387 -701
rect 397 -703 411 -701
rect 441 -703 444 -701
rect 514 -701 523 -699
rect 543 -701 555 -699
rect 580 -701 583 -699
rect 642 -693 651 -691
rect 671 -693 683 -691
rect 723 -693 726 -691
rect 606 -703 608 -700
rect 748 -699 750 -683
rect 851 -689 862 -687
rect 982 -689 994 -687
rect 1004 -689 1007 -687
rect 851 -697 862 -695
rect 982 -697 994 -695
rect 1004 -697 1007 -695
rect 642 -701 651 -699
rect 671 -701 683 -699
rect 723 -701 726 -699
rect 1037 -701 1039 -685
rect 851 -705 862 -703
rect 982 -705 994 -703
rect 1004 -705 1007 -703
rect 377 -711 387 -709
rect 397 -711 411 -709
rect 441 -711 444 -709
rect 152 -717 164 -715
rect 184 -717 200 -715
rect 220 -717 223 -715
rect 473 -712 475 -709
rect 748 -712 750 -709
rect 851 -713 862 -711
rect 982 -713 994 -711
rect 1004 -713 1007 -711
rect 1037 -714 1039 -711
rect 152 -725 164 -723
rect 184 -725 200 -723
rect 220 -725 223 -723
rect 136 -747 138 -744
rect 49 -775 58 -773
rect 78 -775 91 -773
rect 111 -775 114 -773
rect 49 -783 58 -781
rect 78 -783 91 -781
rect 111 -783 114 -781
rect 136 -783 138 -767
rect 136 -796 138 -793
<< polycontact >>
rect 398 225 402 229
rect 398 217 402 221
rect 307 191 311 195
rect 307 183 311 187
rect 494 191 498 195
rect 494 183 498 187
rect 398 169 402 173
rect 398 161 402 165
rect 147 137 151 141
rect 147 129 151 133
rect 56 103 60 107
rect 56 95 60 99
rect 243 103 247 107
rect 243 95 247 99
rect 147 81 151 85
rect 353 84 357 88
rect 147 73 151 77
rect 353 76 357 80
rect 440 80 444 84
rect 471 83 475 87
rect 471 75 475 79
rect 568 80 572 84
rect 44 23 48 27
rect 44 15 48 19
rect 131 19 135 23
rect 276 -2 280 2
rect 276 -10 280 -6
rect 363 -6 367 -2
rect 400 1 404 5
rect 400 -7 404 -3
rect 400 -15 404 -11
rect 516 -13 520 -9
rect 146 -43 150 -39
rect 146 -51 150 -47
rect 55 -77 59 -73
rect 55 -85 59 -81
rect 242 -77 246 -73
rect 242 -85 246 -81
rect 359 -84 363 -80
rect 146 -99 150 -95
rect 359 -92 363 -88
rect 146 -107 150 -103
rect 359 -100 363 -96
rect 437 -92 441 -88
rect 455 -99 459 -95
rect 637 -130 641 -126
rect 637 -138 641 -134
rect 43 -157 47 -153
rect 43 -165 47 -161
rect 130 -161 134 -157
rect 278 -170 282 -166
rect 546 -164 550 -160
rect 278 -178 282 -174
rect 546 -172 550 -168
rect 733 -164 737 -160
rect 733 -172 737 -168
rect 637 -186 641 -182
rect 637 -194 641 -190
rect 187 -204 191 -200
rect 187 -212 191 -208
rect 374 -204 378 -200
rect 374 -212 378 -208
rect 278 -226 282 -222
rect 278 -234 282 -230
rect 533 -268 537 -264
rect 533 -276 537 -272
rect 620 -272 624 -268
rect 146 -297 150 -293
rect 146 -305 150 -301
rect 364 -319 368 -315
rect 55 -331 59 -327
rect 55 -339 59 -335
rect 242 -331 246 -327
rect 364 -327 368 -323
rect 533 -321 537 -317
rect 242 -339 246 -335
rect 364 -335 368 -331
rect 364 -343 368 -339
rect 452 -335 456 -331
rect 470 -337 474 -333
rect 533 -329 537 -325
rect 680 -305 684 -301
rect 680 -313 684 -309
rect 680 -321 684 -317
rect 533 -337 537 -333
rect 629 -336 633 -332
rect 146 -353 150 -349
rect 680 -329 684 -325
rect 817 -325 821 -321
rect 146 -361 150 -357
rect 710 -389 714 -385
rect 779 -388 783 -384
rect 710 -397 714 -393
rect 797 -393 801 -389
rect 43 -411 47 -407
rect 43 -419 47 -415
rect 130 -415 134 -411
rect 292 -432 296 -428
rect 292 -440 296 -436
rect 428 -430 432 -426
rect 292 -448 296 -444
rect 292 -456 296 -452
rect 365 -448 369 -444
rect 384 -449 388 -445
rect 428 -438 432 -434
rect 574 -433 578 -429
rect 428 -446 432 -442
rect 292 -464 296 -460
rect 373 -462 377 -458
rect 428 -454 432 -450
rect 516 -446 520 -442
rect 534 -448 538 -444
rect 574 -441 578 -437
rect 574 -449 578 -445
rect 652 -449 656 -445
rect 670 -448 674 -444
rect 720 -453 724 -449
rect 720 -461 724 -457
rect 720 -469 724 -465
rect 147 -479 151 -475
rect 720 -477 724 -473
rect 875 -469 879 -465
rect 147 -487 151 -483
rect 720 -485 724 -481
rect 56 -513 60 -509
rect 56 -521 60 -517
rect 243 -513 247 -509
rect 243 -521 247 -517
rect 147 -535 151 -531
rect 147 -543 151 -539
rect 470 -548 474 -544
rect 470 -556 474 -552
rect 1095 -551 1099 -547
rect 1095 -559 1099 -555
rect 379 -582 383 -578
rect 44 -593 48 -589
rect 44 -601 48 -597
rect 131 -597 135 -593
rect 379 -590 383 -586
rect 566 -582 570 -578
rect 566 -590 570 -586
rect 470 -604 474 -600
rect 691 -601 695 -597
rect 470 -612 474 -608
rect 691 -609 695 -605
rect 837 -589 841 -585
rect 837 -597 841 -593
rect 924 -593 928 -589
rect 1004 -585 1008 -581
rect 1004 -593 1008 -589
rect 1191 -585 1195 -581
rect 691 -617 695 -613
rect 787 -616 791 -612
rect 1191 -593 1195 -589
rect 1095 -607 1099 -603
rect 1095 -615 1099 -611
rect 148 -662 152 -658
rect 148 -670 152 -666
rect 373 -672 377 -668
rect 373 -680 377 -676
rect 373 -688 377 -684
rect 510 -670 514 -666
rect 510 -678 514 -674
rect 57 -696 61 -692
rect 57 -704 61 -700
rect 244 -696 248 -692
rect 244 -704 248 -700
rect 373 -696 377 -692
rect 444 -688 448 -684
rect 373 -704 377 -700
rect 444 -697 448 -693
rect 469 -696 473 -692
rect 510 -686 514 -682
rect 510 -694 514 -690
rect 583 -686 587 -682
rect 602 -687 606 -683
rect 638 -678 642 -674
rect 638 -686 642 -682
rect 847 -674 851 -670
rect 847 -682 851 -678
rect 148 -718 152 -714
rect 373 -712 377 -708
rect 444 -705 448 -701
rect 510 -702 514 -698
rect 592 -697 596 -693
rect 638 -694 642 -690
rect 638 -702 642 -698
rect 726 -694 730 -690
rect 744 -696 748 -692
rect 847 -690 851 -686
rect 847 -698 851 -694
rect 847 -706 851 -702
rect 1033 -698 1037 -694
rect 847 -714 851 -710
rect 148 -726 152 -722
rect 45 -776 49 -772
rect 45 -784 49 -780
rect 132 -780 136 -776
<< metal1 >>
rect 291 247 504 251
rect 442 236 485 240
rect 405 229 414 233
rect 303 225 398 229
rect 303 195 307 225
rect 394 206 398 221
rect 405 217 408 229
rect 442 225 446 236
rect 470 229 473 233
rect 434 221 446 225
rect 442 217 446 221
rect 351 202 398 206
rect 314 195 323 199
rect 271 191 307 195
rect 271 183 276 191
rect -1 178 276 183
rect 40 159 253 163
rect 191 148 234 152
rect 154 141 163 145
rect 52 137 147 141
rect 52 107 56 137
rect 143 118 147 133
rect 154 129 157 141
rect 191 137 195 148
rect 219 141 222 145
rect 183 133 195 137
rect 191 129 195 133
rect 100 114 147 118
rect 63 107 72 111
rect -1 103 56 107
rect -1 95 12 99
rect 29 27 33 103
rect 45 95 56 99
rect 63 95 66 107
rect 100 103 104 114
rect 128 107 132 111
rect 92 99 104 103
rect 100 95 104 99
rect 52 77 56 95
rect 63 91 72 95
rect 100 91 108 95
rect 143 81 147 114
rect 154 125 163 129
rect 191 125 199 129
rect 154 116 158 125
rect 154 112 203 116
rect 154 89 158 112
rect 230 107 234 148
rect 249 116 253 159
rect 272 143 276 178
rect 288 183 307 187
rect 314 183 317 195
rect 351 191 355 202
rect 379 195 383 199
rect 343 187 355 191
rect 351 183 355 187
rect 288 169 292 183
rect 303 165 307 183
rect 314 179 323 183
rect 351 179 359 183
rect 394 169 398 202
rect 405 213 414 217
rect 442 213 450 217
rect 405 204 409 213
rect 405 200 454 204
rect 405 177 409 200
rect 481 195 485 236
rect 500 204 504 247
rect 538 203 615 207
rect 501 195 510 199
rect 481 191 494 195
rect 481 184 494 187
rect 442 183 494 184
rect 501 183 504 195
rect 538 191 542 203
rect 566 195 570 199
rect 530 187 542 191
rect 538 183 542 187
rect 442 180 485 183
rect 405 173 414 177
rect 303 161 398 165
rect 405 161 408 173
rect 442 169 446 180
rect 501 179 510 183
rect 538 179 546 183
rect 470 173 480 177
rect 434 165 446 169
rect 442 161 446 165
rect 405 157 414 161
rect 442 157 450 161
rect 476 154 480 173
rect 570 154 574 195
rect 291 150 574 154
rect 272 139 346 143
rect 333 119 337 121
rect 287 115 337 119
rect 250 107 259 111
rect 230 103 243 107
rect 230 96 243 99
rect 191 95 243 96
rect 250 95 253 107
rect 287 103 291 115
rect 315 107 319 111
rect 279 99 291 103
rect 287 95 291 99
rect 191 92 234 95
rect 154 85 163 89
rect 52 73 147 77
rect 154 73 157 85
rect 191 81 195 92
rect 250 91 259 95
rect 287 91 295 95
rect 219 85 229 89
rect 183 77 195 81
rect 191 73 195 77
rect 154 69 163 73
rect 191 69 199 73
rect 225 66 229 85
rect 319 66 323 107
rect 333 80 337 115
rect 342 98 346 139
rect 349 116 443 119
rect 467 116 585 119
rect 342 88 346 93
rect 360 92 363 116
rect 439 113 443 116
rect 392 95 432 99
rect 392 92 396 95
rect 360 88 366 92
rect 392 88 399 92
rect 342 84 353 88
rect 333 76 353 80
rect 360 76 363 88
rect 392 84 396 88
rect 428 84 432 95
rect 447 84 451 93
rect 454 84 471 87
rect 386 80 396 84
rect 428 80 440 84
rect 447 83 471 84
rect 447 80 457 83
rect 447 77 451 80
rect 333 72 337 76
rect 360 72 366 76
rect 419 72 425 76
rect 40 62 323 66
rect 422 64 425 72
rect 467 75 471 79
rect 478 75 481 116
rect 567 113 571 116
rect 530 94 558 97
rect 530 91 533 94
rect 524 87 533 91
rect 546 87 552 91
rect 530 83 533 87
rect 530 79 536 83
rect 549 75 552 87
rect 555 84 558 94
rect 575 84 579 93
rect 555 80 568 84
rect 575 80 590 84
rect 575 77 579 80
rect 456 71 471 75
rect 478 71 484 75
rect 546 71 552 75
rect 439 64 443 67
rect 349 61 443 64
rect 40 55 134 58
rect 51 31 54 55
rect 130 52 134 55
rect 83 34 123 38
rect 83 31 87 34
rect 51 27 57 31
rect 83 27 90 31
rect 29 23 44 27
rect 21 15 44 19
rect 51 15 54 27
rect 83 23 87 27
rect 119 23 123 34
rect 138 23 142 32
rect 151 47 444 51
rect 456 51 460 71
rect 549 64 552 71
rect 567 64 571 67
rect 467 61 579 64
rect 449 47 460 51
rect 151 23 155 47
rect 586 34 590 80
rect 272 30 366 33
rect 77 19 87 23
rect 119 19 131 23
rect 138 19 262 23
rect 138 16 142 19
rect 51 11 57 15
rect 110 11 116 15
rect 113 3 116 11
rect 130 3 134 6
rect 40 0 134 3
rect 258 2 262 19
rect 283 6 286 30
rect 362 27 366 30
rect 542 30 590 34
rect 315 9 355 13
rect 315 6 319 9
rect 283 2 289 6
rect 315 2 322 6
rect 258 -2 276 2
rect 262 -10 276 -6
rect 283 -10 286 2
rect 315 -2 319 2
rect 351 -2 355 9
rect 396 23 533 26
rect 370 -2 374 7
rect 381 1 400 5
rect 381 -2 385 1
rect 309 -6 319 -2
rect 351 -6 363 -2
rect 370 -6 385 -2
rect 370 -9 374 -6
rect 388 -7 400 -3
rect 388 -9 392 -7
rect 39 -21 252 -17
rect 190 -32 233 -28
rect 153 -39 162 -35
rect 51 -43 146 -39
rect 51 -73 55 -43
rect 142 -62 146 -47
rect 153 -51 156 -39
rect 190 -43 194 -32
rect 218 -39 221 -35
rect 182 -47 194 -43
rect 190 -51 194 -47
rect 99 -66 146 -62
rect 62 -73 71 -69
rect -2 -77 55 -73
rect -2 -85 11 -81
rect 28 -153 32 -77
rect 44 -85 55 -81
rect 62 -85 65 -73
rect 99 -77 103 -66
rect 127 -73 131 -69
rect 91 -81 103 -77
rect 99 -85 103 -81
rect 51 -103 55 -85
rect 62 -89 71 -85
rect 99 -89 107 -85
rect 142 -99 146 -66
rect 153 -55 162 -51
rect 190 -55 198 -51
rect 153 -64 157 -55
rect 153 -68 202 -64
rect 153 -91 157 -68
rect 229 -73 233 -32
rect 248 -64 252 -21
rect 262 -35 266 -10
rect 283 -14 289 -10
rect 342 -14 348 -10
rect 345 -22 348 -14
rect 382 -13 392 -9
rect 362 -22 366 -19
rect 272 -25 366 -22
rect 262 -39 336 -35
rect 332 -61 336 -39
rect 382 -52 386 -13
rect 396 -42 400 -11
rect 407 -15 410 23
rect 515 20 519 23
rect 479 12 509 15
rect 479 9 482 12
rect 473 5 485 9
rect 479 -7 482 5
rect 498 1 501 9
rect 495 -3 501 1
rect 479 -11 485 -7
rect 498 -15 501 -3
rect 506 -9 509 12
rect 523 -9 527 0
rect 506 -13 516 -9
rect 523 -13 531 -9
rect 407 -19 413 -15
rect 495 -19 501 -15
rect 523 -16 527 -13
rect 407 -25 410 -19
rect 498 -29 501 -19
rect 515 -29 519 -26
rect 424 -32 527 -29
rect 396 -46 491 -42
rect 382 -56 479 -52
rect 286 -65 341 -61
rect 355 -63 472 -60
rect 249 -73 258 -69
rect 229 -77 242 -73
rect 229 -84 242 -81
rect 190 -85 242 -84
rect 249 -85 252 -73
rect 286 -77 290 -65
rect 314 -73 318 -69
rect 278 -81 290 -77
rect 286 -85 290 -81
rect 190 -88 233 -85
rect 153 -95 162 -91
rect 51 -107 146 -103
rect 153 -107 156 -95
rect 190 -99 194 -88
rect 249 -89 258 -85
rect 286 -89 294 -85
rect 218 -95 228 -91
rect 182 -103 194 -99
rect 190 -107 194 -103
rect 153 -111 162 -107
rect 190 -111 198 -107
rect 224 -114 228 -95
rect 286 -102 290 -89
rect 318 -114 322 -73
rect 337 -80 341 -65
rect 337 -84 359 -80
rect 366 -84 369 -63
rect 454 -66 458 -63
rect 398 -73 448 -70
rect 398 -76 401 -73
rect 392 -80 404 -76
rect 329 -88 333 -87
rect 366 -88 372 -84
rect 329 -92 359 -88
rect 347 -100 359 -96
rect 366 -100 369 -88
rect 397 -92 401 -80
rect 392 -96 401 -92
rect 445 -95 448 -73
rect 462 -95 466 -86
rect 475 -95 479 -56
rect 445 -99 455 -95
rect 462 -99 479 -95
rect 366 -104 372 -100
rect 434 -104 440 -100
rect 462 -102 466 -99
rect 39 -118 322 -114
rect 437 -115 440 -104
rect 454 -115 458 -112
rect 355 -118 466 -115
rect 39 -125 133 -122
rect 50 -149 53 -125
rect 129 -128 133 -125
rect 487 -127 491 -46
rect 542 -48 546 30
rect 82 -146 122 -142
rect 82 -149 86 -146
rect 50 -153 56 -149
rect 82 -153 89 -149
rect 28 -157 43 -153
rect 20 -165 43 -161
rect 50 -165 53 -153
rect 82 -157 86 -153
rect 118 -157 122 -146
rect 137 -157 141 -148
rect 150 -131 491 -127
rect 150 -157 154 -131
rect 171 -148 384 -144
rect 76 -161 86 -157
rect 118 -161 130 -157
rect 137 -161 154 -157
rect 322 -159 365 -155
rect 137 -164 141 -161
rect 50 -169 56 -165
rect 109 -169 115 -165
rect 112 -177 115 -169
rect 285 -166 294 -162
rect 183 -170 278 -166
rect 129 -177 133 -174
rect 39 -180 133 -177
rect 183 -200 187 -170
rect 274 -189 278 -174
rect 285 -178 288 -166
rect 322 -170 326 -159
rect 350 -166 353 -162
rect 314 -174 326 -170
rect 322 -178 326 -174
rect 231 -193 278 -189
rect 194 -200 203 -196
rect 165 -204 187 -200
rect 165 -212 187 -208
rect 194 -212 197 -200
rect 231 -204 235 -193
rect 259 -200 263 -196
rect 223 -208 235 -204
rect 231 -212 235 -208
rect 165 -255 168 -212
rect 183 -230 187 -212
rect 194 -216 203 -212
rect 231 -216 239 -212
rect 274 -226 278 -193
rect 285 -182 294 -178
rect 322 -182 330 -178
rect 285 -191 289 -182
rect 285 -195 334 -191
rect 285 -218 289 -195
rect 361 -200 365 -159
rect 380 -191 384 -148
rect 418 -192 472 -188
rect 381 -200 390 -196
rect 361 -204 374 -200
rect 361 -211 374 -208
rect 322 -212 374 -211
rect 381 -212 384 -200
rect 418 -204 422 -192
rect 446 -200 450 -196
rect 410 -208 422 -204
rect 418 -212 422 -208
rect 322 -215 365 -212
rect 285 -222 294 -218
rect 183 -234 278 -230
rect 285 -234 288 -222
rect 322 -226 326 -215
rect 381 -216 390 -212
rect 418 -216 426 -212
rect 350 -222 360 -218
rect 314 -230 326 -226
rect 322 -234 326 -230
rect 285 -238 294 -234
rect 322 -238 330 -234
rect 356 -241 360 -222
rect 450 -241 454 -200
rect 171 -245 454 -241
rect 468 -242 472 -192
rect 487 -235 491 -131
rect 500 -52 546 -48
rect 500 -255 504 -52
rect 611 -84 615 203
rect 611 -88 769 -84
rect 530 -108 743 -104
rect 681 -119 724 -115
rect 644 -126 653 -122
rect 542 -130 637 -126
rect 542 -160 546 -130
rect 633 -149 637 -134
rect 644 -138 647 -126
rect 681 -130 685 -119
rect 709 -126 712 -122
rect 673 -134 685 -130
rect 681 -138 685 -134
rect 590 -153 637 -149
rect 553 -160 562 -156
rect 534 -163 546 -160
rect 530 -164 546 -163
rect 165 -259 504 -255
rect 516 -172 546 -168
rect 553 -172 556 -160
rect 590 -164 594 -153
rect 618 -160 622 -156
rect 582 -168 594 -164
rect 590 -172 594 -168
rect 340 -267 367 -264
rect 39 -275 252 -271
rect 190 -286 233 -282
rect 153 -293 162 -289
rect 51 -297 146 -293
rect 51 -327 55 -297
rect 142 -316 146 -301
rect 153 -305 156 -293
rect 190 -297 194 -286
rect 218 -293 221 -289
rect 182 -301 194 -297
rect 190 -305 194 -301
rect 99 -320 146 -316
rect 62 -327 71 -323
rect -2 -331 55 -327
rect -2 -339 11 -335
rect 28 -407 32 -331
rect 44 -339 55 -335
rect 62 -339 65 -327
rect 99 -331 103 -320
rect 127 -327 131 -323
rect 91 -335 103 -331
rect 99 -339 103 -335
rect 51 -357 55 -339
rect 62 -343 71 -339
rect 99 -343 107 -339
rect 142 -353 146 -320
rect 153 -309 162 -305
rect 190 -309 198 -305
rect 153 -318 157 -309
rect 153 -322 202 -318
rect 153 -345 157 -322
rect 229 -327 233 -286
rect 248 -318 252 -275
rect 340 -287 343 -267
rect 469 -278 472 -268
rect 516 -272 520 -172
rect 542 -190 546 -172
rect 553 -176 562 -172
rect 590 -176 598 -172
rect 633 -186 637 -153
rect 644 -142 653 -138
rect 681 -142 689 -138
rect 644 -151 648 -142
rect 644 -155 693 -151
rect 644 -178 648 -155
rect 720 -160 724 -119
rect 739 -151 743 -108
rect 765 -126 769 -88
rect 765 -130 908 -126
rect 777 -152 892 -148
rect 740 -160 749 -156
rect 720 -164 733 -160
rect 720 -171 733 -168
rect 681 -172 733 -171
rect 740 -172 743 -160
rect 777 -164 781 -152
rect 805 -160 809 -156
rect 769 -168 781 -164
rect 777 -172 781 -168
rect 681 -175 724 -172
rect 644 -182 653 -178
rect 542 -194 637 -190
rect 644 -194 647 -182
rect 681 -186 685 -175
rect 740 -176 749 -172
rect 777 -176 785 -172
rect 709 -182 719 -178
rect 673 -190 685 -186
rect 681 -194 685 -190
rect 644 -198 653 -194
rect 681 -198 689 -194
rect 715 -201 719 -182
rect 809 -201 813 -160
rect 530 -205 813 -201
rect 529 -236 623 -233
rect 529 -268 533 -254
rect 540 -260 543 -236
rect 619 -239 623 -236
rect 572 -257 612 -253
rect 572 -260 576 -257
rect 540 -264 546 -260
rect 572 -264 579 -260
rect 516 -276 533 -272
rect 540 -276 543 -264
rect 572 -268 576 -264
rect 608 -268 612 -257
rect 627 -268 631 -259
rect 566 -272 576 -268
rect 608 -272 620 -268
rect 627 -272 668 -268
rect 627 -275 631 -272
rect 469 -281 494 -278
rect 516 -287 520 -276
rect 540 -280 546 -276
rect 599 -280 605 -276
rect 349 -291 520 -287
rect 602 -288 605 -280
rect 619 -288 623 -285
rect 529 -291 623 -288
rect 349 -295 353 -291
rect 329 -299 353 -295
rect 329 -315 333 -299
rect 360 -301 487 -298
rect 529 -300 646 -297
rect 353 -306 364 -304
rect 353 -308 360 -306
rect 371 -311 374 -301
rect 469 -304 473 -301
rect 403 -308 463 -305
rect 403 -311 406 -308
rect 286 -319 333 -315
rect 344 -318 356 -314
rect 249 -327 258 -323
rect 229 -331 242 -327
rect 229 -338 242 -335
rect 190 -339 242 -338
rect 249 -339 252 -327
rect 286 -331 290 -319
rect 314 -327 318 -323
rect 278 -335 290 -331
rect 286 -339 290 -335
rect 190 -342 233 -339
rect 153 -349 162 -345
rect 51 -361 146 -357
rect 153 -361 156 -349
rect 190 -353 194 -342
rect 249 -343 258 -339
rect 286 -343 294 -339
rect 218 -349 228 -345
rect 182 -357 194 -353
rect 190 -361 194 -357
rect 153 -365 162 -361
rect 190 -365 198 -361
rect 224 -368 228 -349
rect 318 -368 322 -327
rect 329 -339 333 -319
rect 352 -319 356 -318
rect 360 -319 364 -311
rect 371 -315 377 -311
rect 402 -315 409 -311
rect 357 -324 364 -323
rect 352 -327 364 -324
rect 371 -327 374 -315
rect 402 -319 406 -315
rect 397 -323 406 -319
rect 371 -331 377 -327
rect 344 -335 364 -331
rect 329 -343 364 -339
rect 371 -343 374 -331
rect 402 -335 406 -323
rect 460 -333 463 -308
rect 525 -312 533 -308
rect 477 -333 481 -324
rect 397 -339 406 -335
rect 460 -337 470 -333
rect 477 -337 496 -333
rect 477 -340 481 -337
rect 329 -363 333 -343
rect 371 -347 377 -343
rect 449 -347 455 -343
rect 371 -350 374 -347
rect 452 -353 455 -347
rect 469 -353 473 -350
rect 492 -352 496 -337
rect 500 -337 503 -316
rect 529 -321 533 -312
rect 540 -321 543 -300
rect 628 -303 632 -300
rect 664 -301 668 -272
rect 676 -288 834 -285
rect 572 -310 622 -307
rect 572 -313 575 -310
rect 566 -317 578 -313
rect 540 -325 546 -321
rect 515 -328 533 -325
rect 510 -329 533 -328
rect 518 -337 533 -333
rect 540 -337 543 -325
rect 571 -329 575 -317
rect 566 -333 575 -329
rect 611 -337 614 -313
rect 619 -332 622 -310
rect 664 -305 680 -301
rect 659 -313 680 -309
rect 636 -332 640 -323
rect 649 -321 680 -317
rect 649 -332 653 -321
rect 619 -336 629 -332
rect 636 -336 653 -332
rect 661 -329 680 -325
rect 687 -329 690 -288
rect 778 -294 810 -291
rect 778 -297 781 -294
rect 773 -301 781 -297
rect 795 -301 801 -297
rect 777 -305 781 -301
rect 777 -309 785 -305
rect 777 -321 781 -309
rect 798 -313 801 -301
rect 795 -317 801 -313
rect 777 -325 785 -321
rect 798 -329 801 -317
rect 807 -321 810 -294
rect 816 -292 820 -288
rect 824 -321 828 -312
rect 807 -325 817 -321
rect 824 -325 840 -321
rect 824 -328 828 -325
rect 500 -340 508 -337
rect 505 -348 508 -340
rect 360 -356 481 -353
rect 518 -364 522 -337
rect 540 -341 546 -337
rect 608 -341 614 -337
rect 636 -339 640 -336
rect 611 -352 614 -341
rect 628 -352 632 -349
rect 529 -355 640 -352
rect 334 -368 522 -364
rect 661 -362 665 -329
rect 687 -333 693 -329
rect 795 -333 801 -329
rect 798 -341 801 -333
rect 816 -341 820 -338
rect 676 -344 828 -341
rect 706 -357 800 -354
rect 661 -366 710 -362
rect 661 -368 665 -366
rect 39 -372 322 -368
rect 534 -372 665 -368
rect 39 -379 133 -376
rect 50 -403 53 -379
rect 129 -382 133 -379
rect 534 -380 538 -372
rect 82 -400 122 -396
rect 82 -403 86 -400
rect 50 -407 56 -403
rect 82 -407 89 -403
rect 28 -411 43 -407
rect 20 -419 43 -415
rect 50 -419 53 -407
rect 82 -411 86 -407
rect 118 -411 122 -400
rect 137 -411 141 -402
rect 149 -384 538 -380
rect 149 -411 153 -384
rect 706 -389 710 -366
rect 717 -381 720 -357
rect 796 -360 800 -357
rect 749 -378 793 -374
rect 749 -381 753 -378
rect 717 -385 723 -381
rect 749 -385 756 -381
rect 509 -392 684 -389
rect 681 -401 684 -392
rect 698 -396 710 -393
rect 717 -397 720 -385
rect 749 -389 753 -385
rect 743 -393 753 -389
rect 789 -389 793 -378
rect 804 -389 808 -380
rect 836 -381 840 -325
rect 852 -367 855 -344
rect 789 -393 797 -389
rect 804 -393 818 -389
rect 804 -396 808 -393
rect 717 -401 723 -397
rect 776 -401 782 -397
rect 681 -404 699 -401
rect 76 -415 86 -411
rect 118 -415 130 -411
rect 137 -415 153 -411
rect 299 -413 401 -410
rect 424 -412 551 -409
rect 570 -412 687 -409
rect 137 -418 141 -415
rect 50 -423 56 -419
rect 109 -423 115 -419
rect 112 -431 115 -423
rect 129 -431 133 -428
rect 39 -434 133 -431
rect 276 -436 280 -430
rect 288 -432 292 -420
rect 299 -432 302 -413
rect 383 -416 387 -413
rect 331 -421 377 -418
rect 331 -424 334 -421
rect 325 -428 337 -424
rect 299 -436 305 -432
rect 276 -440 292 -436
rect 266 -444 270 -441
rect 266 -448 292 -444
rect 299 -448 302 -436
rect 330 -440 334 -428
rect 325 -444 334 -440
rect 299 -452 305 -448
rect 40 -457 253 -453
rect 257 -456 292 -452
rect 191 -468 234 -464
rect 154 -475 163 -471
rect 52 -479 147 -475
rect 52 -509 56 -479
rect 143 -498 147 -483
rect 154 -487 157 -475
rect 191 -479 195 -468
rect 219 -475 222 -471
rect 183 -483 195 -479
rect 191 -487 195 -483
rect 100 -502 147 -498
rect 63 -509 72 -505
rect -1 -513 56 -509
rect -1 -521 12 -517
rect 29 -589 33 -513
rect 45 -521 56 -517
rect 63 -521 66 -509
rect 100 -513 104 -502
rect 128 -509 132 -505
rect 92 -517 104 -513
rect 100 -521 104 -517
rect 52 -539 56 -521
rect 63 -525 72 -521
rect 100 -525 108 -521
rect 143 -535 147 -502
rect 154 -491 163 -487
rect 191 -491 199 -487
rect 154 -500 158 -491
rect 154 -504 203 -500
rect 154 -527 158 -504
rect 230 -509 234 -468
rect 249 -500 253 -457
rect 268 -488 272 -456
rect 280 -464 292 -460
rect 299 -464 302 -452
rect 330 -456 334 -444
rect 374 -445 377 -421
rect 425 -422 428 -417
rect 424 -430 428 -422
rect 435 -422 438 -412
rect 533 -415 537 -412
rect 467 -419 527 -416
rect 467 -422 470 -419
rect 435 -426 441 -422
rect 466 -426 473 -422
rect 391 -445 395 -436
rect 402 -435 428 -434
rect 407 -438 428 -435
rect 435 -438 438 -426
rect 466 -430 470 -426
rect 461 -434 470 -430
rect 435 -442 441 -438
rect 411 -445 428 -442
rect 374 -449 384 -445
rect 391 -449 406 -445
rect 391 -452 395 -449
rect 325 -460 334 -456
rect 280 -491 284 -464
rect 299 -468 305 -464
rect 362 -465 365 -464
rect 362 -468 368 -465
rect 365 -474 368 -468
rect 383 -474 387 -462
rect 288 -477 387 -474
rect 402 -480 406 -449
rect 416 -446 428 -445
rect 424 -462 428 -450
rect 435 -454 438 -442
rect 466 -446 470 -434
rect 524 -444 527 -419
rect 566 -423 574 -419
rect 570 -433 574 -423
rect 581 -433 584 -412
rect 669 -415 673 -412
rect 613 -422 663 -419
rect 613 -425 616 -422
rect 607 -429 619 -425
rect 541 -444 545 -435
rect 581 -437 587 -433
rect 557 -441 574 -437
rect 461 -450 470 -446
rect 524 -448 534 -444
rect 541 -447 559 -444
rect 541 -448 546 -447
rect 551 -448 559 -447
rect 541 -451 545 -448
rect 435 -458 441 -454
rect 513 -455 516 -454
rect 513 -458 519 -455
rect 435 -461 438 -458
rect 516 -464 519 -458
rect 533 -464 537 -461
rect 439 -467 545 -464
rect 555 -478 559 -448
rect 567 -449 574 -445
rect 581 -449 584 -437
rect 612 -441 616 -429
rect 607 -445 616 -441
rect 660 -444 663 -422
rect 696 -420 699 -404
rect 779 -409 782 -401
rect 796 -409 800 -406
rect 706 -412 800 -409
rect 814 -415 818 -393
rect 888 -390 892 -152
rect 904 -375 908 -130
rect 904 -379 935 -375
rect 888 -394 919 -390
rect 829 -397 877 -394
rect 874 -409 877 -397
rect 874 -412 892 -409
rect 709 -419 818 -415
rect 677 -444 681 -435
rect 709 -442 713 -419
rect 822 -425 907 -422
rect 716 -433 892 -430
rect 660 -448 670 -444
rect 677 -448 686 -444
rect 709 -446 720 -442
rect 567 -458 571 -449
rect 581 -453 587 -449
rect 618 -453 619 -449
rect 677 -451 681 -448
rect 618 -464 621 -453
rect 716 -453 720 -446
rect 709 -461 720 -457
rect 669 -464 673 -461
rect 597 -467 681 -464
rect 708 -469 720 -465
rect 580 -476 679 -472
rect 333 -486 364 -482
rect 402 -484 459 -480
rect 280 -495 291 -491
rect 287 -497 291 -495
rect 333 -497 337 -486
rect 580 -490 584 -476
rect 287 -501 337 -497
rect 345 -494 584 -490
rect 250 -509 259 -505
rect 230 -513 243 -509
rect 230 -520 243 -517
rect 191 -521 243 -520
rect 250 -521 253 -509
rect 287 -513 291 -501
rect 315 -509 319 -505
rect 345 -505 349 -494
rect 331 -509 349 -505
rect 279 -517 291 -513
rect 287 -521 291 -517
rect 191 -524 234 -521
rect 154 -531 163 -527
rect 52 -543 147 -539
rect 154 -543 157 -531
rect 191 -535 195 -524
rect 250 -525 259 -521
rect 287 -525 295 -521
rect 219 -531 229 -527
rect 183 -539 195 -535
rect 191 -543 195 -539
rect 154 -547 163 -543
rect 191 -547 199 -543
rect 225 -550 229 -531
rect 287 -535 291 -525
rect 260 -541 286 -537
rect 319 -550 323 -509
rect 40 -554 323 -550
rect 331 -558 335 -509
rect 363 -526 576 -522
rect 514 -537 557 -533
rect 477 -544 486 -540
rect 40 -561 134 -558
rect 51 -585 54 -561
rect 130 -564 134 -561
rect 151 -562 335 -558
rect 375 -548 470 -544
rect 83 -582 123 -578
rect 83 -585 87 -582
rect 51 -589 57 -585
rect 83 -589 90 -585
rect 29 -593 44 -589
rect 21 -601 44 -597
rect 51 -601 54 -589
rect 83 -593 87 -589
rect 119 -593 123 -582
rect 138 -593 142 -584
rect 151 -593 155 -562
rect 77 -597 87 -593
rect 119 -597 131 -593
rect 138 -597 155 -593
rect 138 -600 142 -597
rect 51 -605 57 -601
rect 110 -605 116 -601
rect 113 -613 116 -605
rect 130 -613 134 -610
rect 40 -616 134 -613
rect 256 -625 259 -570
rect 268 -609 272 -572
rect 315 -574 367 -570
rect 363 -578 367 -574
rect 375 -578 379 -548
rect 466 -567 470 -552
rect 477 -556 480 -544
rect 514 -548 518 -537
rect 542 -544 545 -540
rect 506 -552 518 -548
rect 514 -556 518 -552
rect 423 -571 470 -567
rect 386 -578 395 -574
rect 363 -582 379 -578
rect 334 -586 339 -585
rect 334 -590 379 -586
rect 386 -590 389 -578
rect 423 -582 427 -571
rect 451 -578 455 -574
rect 415 -586 427 -582
rect 423 -590 427 -586
rect 283 -598 346 -595
rect 268 -612 337 -609
rect 268 -613 272 -612
rect 256 -628 325 -625
rect 41 -640 254 -636
rect 192 -651 235 -647
rect 155 -658 164 -654
rect 53 -662 148 -658
rect 53 -692 57 -662
rect 144 -681 148 -666
rect 155 -670 158 -658
rect 192 -662 196 -651
rect 220 -658 223 -654
rect 184 -666 196 -662
rect 192 -670 196 -666
rect 101 -685 148 -681
rect 64 -692 73 -688
rect 0 -696 57 -692
rect 0 -704 13 -700
rect 30 -772 34 -696
rect 46 -704 57 -700
rect 64 -704 67 -692
rect 101 -696 105 -685
rect 129 -692 133 -688
rect 93 -700 105 -696
rect 101 -704 105 -700
rect 53 -722 57 -704
rect 64 -708 73 -704
rect 101 -708 109 -704
rect 144 -718 148 -685
rect 155 -674 164 -670
rect 192 -674 200 -670
rect 155 -683 159 -674
rect 155 -687 204 -683
rect 155 -710 159 -687
rect 231 -692 235 -651
rect 250 -683 254 -640
rect 322 -679 325 -628
rect 334 -663 337 -612
rect 322 -682 331 -679
rect 251 -692 260 -688
rect 231 -696 244 -692
rect 231 -703 244 -700
rect 192 -704 244 -703
rect 251 -704 254 -692
rect 288 -696 292 -684
rect 316 -692 320 -688
rect 280 -700 292 -696
rect 288 -704 292 -700
rect 192 -707 235 -704
rect 155 -714 164 -710
rect 53 -726 148 -722
rect 155 -726 158 -714
rect 192 -718 196 -707
rect 251 -708 260 -704
rect 288 -708 296 -704
rect 220 -714 230 -710
rect 184 -722 196 -718
rect 192 -726 196 -722
rect 155 -730 164 -726
rect 192 -730 200 -726
rect 226 -733 230 -714
rect 288 -718 292 -708
rect 288 -722 302 -718
rect 320 -733 324 -692
rect 328 -700 331 -682
rect 343 -684 346 -598
rect 375 -608 379 -590
rect 386 -594 395 -590
rect 423 -594 431 -590
rect 466 -604 470 -571
rect 477 -560 486 -556
rect 514 -560 522 -556
rect 477 -569 481 -560
rect 477 -573 526 -569
rect 477 -596 481 -573
rect 553 -578 557 -537
rect 572 -569 576 -526
rect 655 -552 659 -476
rect 675 -496 679 -476
rect 707 -477 720 -473
rect 707 -486 711 -477
rect 700 -490 711 -486
rect 716 -496 720 -481
rect 727 -485 730 -433
rect 874 -436 878 -433
rect 839 -442 868 -439
rect 839 -445 842 -442
rect 833 -449 845 -445
rect 838 -461 842 -449
rect 858 -453 861 -445
rect 855 -457 861 -453
rect 838 -465 845 -461
rect 838 -477 842 -465
rect 858 -469 861 -457
rect 865 -465 868 -442
rect 882 -465 886 -456
rect 865 -469 875 -465
rect 882 -469 893 -465
rect 855 -473 861 -469
rect 882 -472 886 -469
rect 838 -481 845 -477
rect 858 -485 861 -473
rect 727 -489 733 -485
rect 855 -486 861 -485
rect 874 -486 878 -482
rect 855 -489 878 -486
rect 727 -495 730 -489
rect 675 -500 720 -496
rect 858 -499 861 -489
rect 739 -502 861 -499
rect 904 -506 907 -425
rect 915 -450 919 -394
rect 931 -437 935 -379
rect 931 -441 963 -437
rect 915 -454 948 -450
rect 944 -496 948 -454
rect 959 -465 963 -441
rect 959 -469 1284 -465
rect 958 -489 1285 -485
rect 944 -500 1285 -496
rect 679 -509 907 -506
rect 948 -509 1285 -505
rect 655 -556 665 -552
rect 610 -570 668 -566
rect 573 -578 582 -574
rect 553 -582 566 -578
rect 553 -589 566 -586
rect 514 -590 566 -589
rect 573 -590 576 -578
rect 610 -582 614 -570
rect 638 -578 642 -574
rect 602 -586 614 -582
rect 610 -590 614 -586
rect 514 -593 557 -590
rect 477 -600 486 -596
rect 375 -612 470 -608
rect 477 -612 480 -600
rect 514 -604 518 -593
rect 573 -594 582 -590
rect 610 -594 618 -590
rect 542 -600 552 -596
rect 506 -608 518 -604
rect 514 -612 518 -608
rect 477 -616 486 -612
rect 514 -616 522 -612
rect 548 -619 552 -600
rect 642 -619 646 -578
rect 679 -597 682 -509
rect 948 -521 952 -509
rect 785 -525 952 -521
rect 785 -566 789 -525
rect 988 -529 1201 -525
rect 1139 -540 1182 -536
rect 833 -557 927 -554
rect 695 -569 789 -566
rect 694 -570 789 -569
rect 687 -580 804 -577
rect 679 -601 691 -597
rect 698 -601 701 -580
rect 786 -583 790 -580
rect 730 -590 780 -587
rect 730 -593 733 -590
rect 724 -597 736 -593
rect 698 -605 704 -601
rect 676 -609 691 -605
rect 363 -623 646 -619
rect 687 -620 691 -613
rect 698 -617 701 -605
rect 729 -609 733 -597
rect 724 -613 733 -609
rect 769 -617 772 -593
rect 777 -612 780 -590
rect 811 -585 815 -557
rect 844 -581 847 -557
rect 923 -560 927 -557
rect 876 -578 916 -574
rect 876 -581 880 -578
rect 844 -585 850 -581
rect 876 -585 883 -581
rect 811 -589 837 -585
rect 814 -594 837 -593
rect 819 -597 837 -594
rect 844 -597 847 -585
rect 876 -589 880 -585
rect 912 -589 916 -578
rect 931 -589 935 -580
rect 988 -581 992 -545
rect 1102 -547 1111 -543
rect 1000 -551 1095 -547
rect 1000 -581 1004 -551
rect 1091 -570 1095 -555
rect 1102 -559 1105 -547
rect 1139 -551 1143 -540
rect 1167 -547 1170 -543
rect 1131 -555 1143 -551
rect 1139 -559 1143 -555
rect 1048 -574 1095 -570
rect 1011 -581 1020 -577
rect 988 -585 1004 -581
rect 870 -593 880 -589
rect 912 -593 924 -589
rect 931 -593 952 -589
rect 931 -596 935 -593
rect 844 -601 850 -597
rect 903 -601 909 -597
rect 794 -612 798 -603
rect 906 -609 909 -601
rect 923 -609 927 -606
rect 833 -612 927 -609
rect 777 -616 787 -612
rect 794 -616 826 -612
rect 667 -623 691 -620
rect 698 -621 704 -617
rect 766 -621 772 -617
rect 794 -619 798 -616
rect 769 -632 772 -621
rect 786 -632 790 -629
rect 710 -635 798 -632
rect 380 -649 472 -645
rect 362 -664 373 -660
rect 369 -672 373 -664
rect 380 -664 384 -649
rect 403 -661 465 -657
rect 403 -664 407 -661
rect 380 -668 387 -664
rect 403 -668 411 -664
rect 359 -676 363 -672
rect 359 -680 373 -676
rect 380 -680 384 -668
rect 403 -672 407 -668
rect 397 -676 407 -672
rect 380 -684 387 -680
rect 343 -688 373 -684
rect 339 -694 373 -692
rect 334 -696 373 -694
rect 380 -696 384 -684
rect 403 -688 407 -676
rect 397 -692 407 -688
rect 461 -692 465 -661
rect 468 -663 472 -649
rect 506 -651 604 -648
rect 507 -661 510 -656
rect 506 -670 510 -661
rect 517 -670 520 -651
rect 601 -654 605 -651
rect 549 -659 598 -656
rect 549 -662 552 -659
rect 543 -666 555 -662
rect 517 -674 523 -670
rect 497 -678 510 -674
rect 380 -700 387 -696
rect 328 -704 373 -700
rect 335 -710 373 -708
rect 340 -712 373 -710
rect 380 -712 384 -700
rect 403 -704 407 -692
rect 461 -696 469 -692
rect 476 -699 480 -683
rect 492 -686 510 -682
rect 517 -686 520 -674
rect 548 -678 552 -666
rect 543 -682 552 -678
rect 492 -687 497 -686
rect 397 -708 407 -704
rect 468 -712 472 -709
rect 380 -716 387 -712
rect 441 -715 472 -712
rect 502 -701 505 -691
rect 517 -690 523 -686
rect 441 -716 444 -715
rect 380 -722 384 -716
rect 41 -737 324 -733
rect 41 -744 135 -741
rect 476 -743 480 -709
rect 511 -710 514 -702
rect 517 -702 520 -690
rect 548 -694 552 -682
rect 595 -683 598 -659
rect 634 -660 761 -657
rect 822 -660 826 -616
rect 948 -618 952 -593
rect 978 -593 1004 -589
rect 1011 -593 1014 -581
rect 1048 -585 1052 -574
rect 1076 -581 1080 -577
rect 1040 -589 1052 -585
rect 1048 -593 1052 -589
rect 1000 -611 1004 -593
rect 1011 -597 1020 -593
rect 1048 -597 1056 -593
rect 1091 -607 1095 -574
rect 1102 -563 1111 -559
rect 1139 -563 1147 -559
rect 1102 -572 1106 -563
rect 1102 -576 1151 -572
rect 1102 -599 1106 -576
rect 1178 -581 1182 -540
rect 1197 -572 1201 -529
rect 1235 -573 1285 -569
rect 1198 -581 1207 -577
rect 1178 -585 1191 -581
rect 1178 -592 1191 -589
rect 1139 -593 1191 -592
rect 1198 -593 1201 -581
rect 1235 -585 1239 -573
rect 1263 -581 1267 -577
rect 1227 -589 1239 -585
rect 1235 -593 1239 -589
rect 1139 -596 1182 -593
rect 1102 -603 1111 -599
rect 1000 -615 1095 -611
rect 1102 -615 1105 -603
rect 1139 -607 1143 -596
rect 1198 -597 1207 -593
rect 1235 -597 1243 -593
rect 1167 -603 1177 -599
rect 1131 -611 1143 -607
rect 1139 -615 1143 -611
rect 842 -622 952 -618
rect 1102 -619 1111 -615
rect 1139 -619 1147 -615
rect 1173 -622 1177 -603
rect 1267 -622 1271 -581
rect 645 -670 648 -660
rect 743 -663 747 -660
rect 822 -663 833 -660
rect 677 -667 737 -664
rect 677 -670 680 -667
rect 595 -687 602 -683
rect 609 -690 613 -674
rect 635 -675 638 -670
rect 645 -674 651 -670
rect 676 -674 683 -670
rect 634 -678 638 -675
rect 623 -684 638 -682
rect 628 -686 638 -684
rect 645 -686 648 -674
rect 676 -678 680 -674
rect 671 -682 680 -678
rect 645 -690 651 -686
rect 543 -698 552 -694
rect 517 -706 523 -702
rect 580 -706 586 -702
rect 583 -712 586 -706
rect 601 -712 605 -700
rect 532 -715 605 -712
rect 634 -692 638 -690
rect 609 -724 613 -700
rect 622 -695 638 -692
rect 622 -696 627 -695
rect 645 -702 648 -690
rect 676 -694 680 -682
rect 734 -692 737 -667
rect 829 -666 833 -663
rect 842 -670 846 -622
rect 988 -626 1271 -622
rect 1277 -582 1286 -578
rect 1277 -632 1281 -582
rect 1057 -636 1281 -632
rect 854 -654 1029 -650
rect 842 -674 847 -670
rect 751 -692 755 -683
rect 768 -682 847 -678
rect 768 -692 772 -682
rect 671 -698 680 -694
rect 734 -696 744 -692
rect 751 -696 772 -692
rect 785 -690 847 -686
rect 751 -699 755 -696
rect 645 -706 651 -702
rect 723 -706 729 -702
rect 645 -709 648 -706
rect 726 -712 729 -706
rect 743 -712 747 -709
rect 634 -715 755 -712
rect 785 -724 789 -690
rect 609 -728 789 -724
rect 797 -698 847 -694
rect 797 -743 801 -698
rect 835 -706 847 -702
rect 843 -716 847 -710
rect 854 -714 858 -654
rect 985 -662 1022 -658
rect 1026 -659 1029 -654
rect 1026 -662 1036 -659
rect 985 -666 989 -662
rect 982 -670 989 -666
rect 1004 -670 1011 -666
rect 985 -674 989 -670
rect 985 -678 994 -674
rect 985 -690 989 -678
rect 1007 -682 1011 -670
rect 1004 -686 1011 -682
rect 985 -694 994 -690
rect 985 -706 989 -694
rect 1007 -698 1011 -686
rect 1018 -694 1022 -662
rect 1032 -665 1036 -662
rect 1040 -694 1044 -685
rect 1057 -694 1061 -636
rect 1018 -698 1033 -694
rect 1040 -698 1061 -694
rect 1004 -702 1011 -698
rect 1040 -701 1044 -698
rect 985 -710 994 -706
rect 1007 -713 1011 -702
rect 1032 -713 1036 -711
rect 1007 -714 1036 -713
rect 52 -768 55 -744
rect 131 -747 135 -744
rect 154 -747 438 -743
rect 476 -747 801 -743
rect 811 -720 847 -716
rect 854 -718 862 -714
rect 1004 -717 1036 -714
rect 1004 -718 1011 -717
rect 84 -765 124 -761
rect 84 -768 88 -765
rect 52 -772 58 -768
rect 84 -772 91 -768
rect 30 -776 45 -772
rect 22 -784 45 -780
rect 52 -784 55 -772
rect 84 -776 88 -772
rect 120 -776 124 -765
rect 139 -776 143 -767
rect 154 -776 158 -747
rect 434 -752 438 -747
rect 811 -752 815 -720
rect 434 -756 815 -752
rect 78 -780 88 -776
rect 120 -780 132 -776
rect 139 -780 158 -776
rect 139 -783 143 -780
rect 52 -788 58 -784
rect 111 -788 117 -784
rect 114 -796 117 -788
rect 131 -796 135 -793
rect 41 -799 135 -796
<< m2contact >>
rect 313 242 318 247
rect 473 228 478 233
rect 313 199 318 204
rect 62 154 67 159
rect 222 140 227 145
rect 62 111 67 116
rect 12 95 17 100
rect 40 95 45 100
rect 132 106 137 111
rect 203 112 208 117
rect 383 194 388 199
rect 287 164 292 169
rect 454 200 459 205
rect 499 199 504 204
rect 570 195 575 200
rect 333 121 338 126
rect 248 111 253 116
rect 319 107 324 112
rect 342 93 347 98
rect 332 66 338 72
rect 21 19 26 24
rect 444 47 449 52
rect 61 -26 66 -21
rect 221 -40 226 -35
rect 61 -69 66 -64
rect 11 -85 16 -80
rect 39 -85 44 -80
rect 131 -74 136 -69
rect 202 -68 207 -63
rect 531 -13 536 -8
rect 247 -69 252 -64
rect 318 -73 323 -68
rect 286 -107 291 -102
rect 328 -87 333 -82
rect 342 -101 347 -96
rect 437 -97 442 -92
rect 20 -161 25 -156
rect 193 -153 198 -148
rect 165 -200 170 -195
rect 353 -167 358 -162
rect 193 -196 198 -191
rect 263 -201 268 -196
rect 334 -195 339 -190
rect 379 -196 384 -191
rect 450 -200 455 -195
rect 487 -240 492 -235
rect 468 -247 473 -242
rect 552 -113 557 -108
rect 529 -163 534 -158
rect 712 -127 717 -122
rect 552 -156 557 -151
rect 622 -161 627 -156
rect 61 -280 66 -275
rect 221 -294 226 -289
rect 61 -323 66 -318
rect 11 -339 16 -334
rect 39 -339 44 -334
rect 131 -328 136 -323
rect 202 -322 207 -317
rect 367 -269 372 -264
rect 468 -268 473 -263
rect 693 -155 698 -150
rect 738 -156 743 -151
rect 809 -160 814 -155
rect 529 -254 534 -249
rect 494 -282 499 -277
rect 339 -292 344 -287
rect 348 -308 353 -303
rect 360 -311 365 -306
rect 247 -323 252 -318
rect 339 -318 344 -313
rect 318 -327 323 -322
rect 352 -324 357 -319
rect 339 -334 344 -329
rect 499 -316 504 -311
rect 520 -312 525 -307
rect 452 -340 457 -335
rect 510 -328 515 -323
rect 653 -314 659 -308
rect 491 -358 497 -352
rect 504 -353 509 -348
rect 329 -368 334 -363
rect 20 -415 25 -410
rect 504 -394 509 -389
rect 693 -397 698 -392
rect 779 -394 785 -388
rect 851 -344 856 -339
rect 851 -372 856 -367
rect 836 -386 841 -381
rect 287 -420 292 -415
rect 276 -430 281 -425
rect 266 -441 271 -436
rect 257 -452 262 -447
rect 62 -462 67 -457
rect 222 -476 227 -471
rect 62 -505 67 -500
rect 12 -521 17 -516
rect 40 -521 45 -516
rect 132 -510 137 -505
rect 203 -504 208 -499
rect 420 -422 425 -417
rect 402 -440 407 -435
rect 365 -453 370 -448
rect 267 -494 273 -488
rect 373 -467 378 -462
rect 411 -450 416 -445
rect 561 -423 566 -418
rect 552 -441 557 -436
rect 516 -451 521 -446
rect 423 -467 428 -462
rect 652 -445 657 -440
rect 824 -399 829 -394
rect 892 -413 897 -408
rect 695 -425 700 -420
rect 817 -427 822 -422
rect 686 -448 691 -443
rect 567 -463 572 -458
rect 704 -461 709 -456
rect 703 -470 708 -465
rect 364 -486 369 -481
rect 459 -484 464 -479
rect 554 -484 560 -478
rect 248 -505 253 -500
rect 319 -509 324 -504
rect 254 -541 260 -535
rect 286 -541 292 -535
rect 385 -531 390 -526
rect 21 -597 26 -592
rect 255 -570 260 -565
rect 267 -572 273 -566
rect 309 -575 315 -569
rect 545 -545 550 -540
rect 385 -574 390 -569
rect 334 -585 339 -580
rect 455 -579 460 -574
rect 278 -600 283 -595
rect 63 -645 68 -640
rect 223 -659 228 -654
rect 63 -688 68 -683
rect 13 -704 18 -699
rect 41 -704 46 -699
rect 133 -693 138 -688
rect 204 -687 209 -682
rect 333 -668 338 -663
rect 249 -688 254 -683
rect 320 -692 325 -687
rect 302 -722 307 -717
rect 526 -573 531 -568
rect 695 -491 700 -486
rect 893 -470 899 -464
rect 953 -490 958 -485
rect 665 -557 671 -551
rect 571 -574 576 -569
rect 668 -570 673 -565
rect 642 -578 647 -573
rect 690 -569 695 -564
rect 1010 -534 1015 -529
rect 987 -545 993 -539
rect 810 -557 816 -551
rect 676 -614 681 -609
rect 814 -599 819 -594
rect 1170 -548 1175 -543
rect 1010 -577 1015 -572
rect 662 -625 667 -620
rect 357 -664 362 -659
rect 354 -677 359 -672
rect 334 -694 339 -689
rect 448 -688 453 -683
rect 502 -661 507 -656
rect 492 -679 497 -674
rect 335 -715 340 -710
rect 448 -697 453 -692
rect 492 -692 497 -687
rect 448 -706 453 -701
rect 505 -694 510 -689
rect 501 -706 506 -701
rect 973 -594 978 -589
rect 1080 -582 1085 -577
rect 1151 -576 1156 -571
rect 1196 -577 1201 -572
rect 1267 -581 1272 -576
rect 583 -691 588 -686
rect 630 -675 635 -670
rect 623 -689 628 -684
rect 592 -702 597 -697
rect 509 -715 514 -710
rect 622 -701 627 -696
rect 637 -707 642 -702
rect 726 -690 731 -685
rect 828 -672 834 -666
rect 827 -709 835 -701
rect 22 -780 27 -775
<< metal2 >>
rect 314 204 317 242
rect 475 221 478 228
rect 475 218 574 221
rect 475 212 478 218
rect 447 209 478 212
rect 447 198 450 209
rect 459 201 499 204
rect 571 200 574 218
rect 388 195 450 198
rect 63 116 66 154
rect 283 148 287 169
rect 283 144 337 148
rect 224 133 227 140
rect 239 133 323 136
rect 224 130 242 133
rect 224 124 227 130
rect 196 121 227 124
rect 196 110 199 121
rect 208 113 248 116
rect 320 112 323 133
rect 333 126 337 144
rect 137 107 199 110
rect 17 95 40 99
rect 21 24 25 95
rect 62 -64 65 -26
rect 223 -47 226 -40
rect 223 -50 322 -47
rect 223 -56 226 -50
rect 195 -59 226 -56
rect 195 -70 198 -59
rect 207 -67 247 -64
rect 319 -68 322 -50
rect 333 -51 337 66
rect 328 -55 337 -51
rect 136 -73 198 -70
rect 16 -85 39 -81
rect 328 -82 332 -55
rect 20 -156 24 -85
rect 343 -96 346 93
rect 445 -38 448 47
rect 536 -11 554 -8
rect 378 -41 448 -38
rect 378 -75 381 -41
rect 551 -57 554 -11
rect 511 -60 554 -57
rect 378 -78 481 -75
rect 442 -97 444 -92
rect 287 -133 290 -107
rect 166 -136 290 -133
rect 166 -184 169 -136
rect 343 -143 346 -101
rect 251 -146 346 -143
rect 155 -187 169 -184
rect 155 -269 158 -187
rect 166 -195 169 -187
rect 194 -191 197 -153
rect 251 -261 254 -146
rect 441 -156 444 -97
rect 441 -159 460 -156
rect 355 -174 358 -167
rect 457 -166 460 -159
rect 457 -169 463 -166
rect 355 -177 454 -174
rect 355 -183 358 -177
rect 327 -186 358 -183
rect 327 -197 330 -186
rect 339 -194 379 -191
rect 451 -195 454 -177
rect 268 -200 330 -197
rect 460 -208 463 -169
rect 457 -211 463 -208
rect 251 -264 352 -261
rect 155 -272 330 -269
rect 62 -318 65 -280
rect 223 -301 226 -294
rect 223 -304 322 -301
rect 223 -310 226 -304
rect 195 -313 226 -310
rect 195 -324 198 -313
rect 207 -321 247 -318
rect 319 -322 322 -304
rect 136 -327 198 -324
rect 327 -330 330 -272
rect 340 -313 343 -292
rect 349 -303 352 -264
rect 457 -265 460 -211
rect 478 -218 481 -78
rect 511 -159 514 -60
rect 553 -151 556 -113
rect 714 -134 717 -127
rect 714 -137 813 -134
rect 714 -143 717 -137
rect 686 -146 717 -143
rect 511 -162 529 -159
rect 686 -157 689 -146
rect 698 -154 738 -151
rect 810 -155 813 -137
rect 627 -160 689 -157
rect 478 -221 684 -218
rect 469 -263 472 -247
rect 372 -268 460 -265
rect 478 -265 481 -221
rect 492 -238 519 -235
rect 516 -241 519 -238
rect 516 -242 532 -241
rect 516 -244 542 -242
rect 529 -245 667 -244
rect 529 -249 532 -245
rect 539 -247 667 -245
rect 478 -268 511 -265
rect 478 -277 481 -268
rect 421 -280 481 -277
rect 327 -333 339 -330
rect 16 -339 39 -335
rect 20 -410 24 -339
rect 336 -345 339 -333
rect 248 -348 346 -345
rect 248 -445 251 -348
rect 330 -386 333 -368
rect 102 -448 251 -445
rect 258 -389 333 -386
rect 258 -447 261 -389
rect 343 -393 346 -348
rect 267 -396 346 -393
rect 267 -436 270 -396
rect 353 -400 356 -324
rect 277 -403 356 -400
rect 277 -425 280 -403
rect 361 -408 364 -311
rect 288 -411 364 -408
rect 288 -415 291 -411
rect 63 -500 66 -462
rect 17 -521 40 -517
rect 21 -592 25 -521
rect 102 -578 105 -448
rect 277 -460 280 -430
rect 111 -463 280 -460
rect 111 -570 114 -463
rect 224 -483 227 -476
rect 257 -479 280 -476
rect 257 -483 260 -479
rect 224 -486 260 -483
rect 277 -483 280 -479
rect 277 -486 323 -483
rect 224 -492 227 -486
rect 196 -495 227 -492
rect 196 -506 199 -495
rect 208 -503 248 -500
rect 137 -509 199 -506
rect 255 -565 259 -541
rect 268 -566 272 -494
rect 320 -504 323 -486
rect 111 -573 235 -570
rect 287 -570 291 -541
rect 102 -581 228 -578
rect 225 -596 228 -581
rect 232 -583 235 -573
rect 287 -574 309 -570
rect 328 -573 331 -411
rect 421 -417 424 -280
rect 495 -311 498 -282
rect 508 -304 511 -268
rect 508 -307 524 -304
rect 495 -315 499 -311
rect 497 -328 510 -325
rect 497 -336 500 -328
rect 457 -339 500 -336
rect 483 -340 487 -339
rect 492 -399 496 -358
rect 505 -389 508 -353
rect 654 -360 658 -314
rect 524 -364 658 -360
rect 664 -351 667 -247
rect 681 -272 684 -221
rect 681 -275 855 -272
rect 852 -339 855 -275
rect 852 -345 855 -344
rect 664 -354 870 -351
rect 524 -399 528 -364
rect 664 -375 667 -354
rect 852 -367 855 -366
rect 562 -378 667 -375
rect 492 -401 497 -399
rect 524 -401 529 -399
rect 492 -405 529 -401
rect 562 -418 565 -378
rect 654 -396 693 -393
rect 403 -449 406 -440
rect 654 -440 657 -396
rect 700 -423 769 -420
rect 766 -434 769 -423
rect 785 -423 788 -388
rect 822 -399 824 -395
rect 822 -407 825 -399
rect 822 -410 833 -407
rect 785 -426 817 -423
rect 830 -434 833 -410
rect 766 -437 833 -434
rect 370 -452 406 -449
rect 412 -464 415 -450
rect 553 -447 556 -441
rect 521 -450 556 -447
rect 687 -458 690 -448
rect 378 -467 415 -464
rect 687 -461 704 -458
rect 424 -471 427 -467
rect 568 -471 571 -463
rect 424 -474 571 -471
rect 424 -481 427 -474
rect 369 -484 427 -481
rect 703 -479 706 -470
rect 580 -480 706 -479
rect 560 -482 706 -480
rect 560 -483 584 -482
rect 460 -498 463 -484
rect 587 -490 695 -487
rect 587 -498 590 -490
rect 460 -501 590 -498
rect 837 -508 840 -386
rect 324 -576 331 -573
rect 335 -511 840 -508
rect 232 -586 310 -583
rect 225 -599 278 -596
rect 307 -606 310 -586
rect 324 -598 327 -576
rect 335 -580 338 -511
rect 852 -526 855 -372
rect 439 -529 855 -526
rect 386 -569 389 -531
rect 324 -601 360 -598
rect 307 -609 352 -606
rect 64 -683 67 -645
rect 225 -666 228 -659
rect 349 -657 352 -609
rect 357 -648 360 -601
rect 439 -633 442 -529
rect 867 -538 870 -354
rect 897 -411 957 -408
rect 899 -469 923 -465
rect 547 -552 550 -545
rect 653 -541 870 -538
rect 919 -540 923 -469
rect 954 -485 957 -411
rect 547 -555 646 -552
rect 547 -561 550 -555
rect 519 -564 550 -561
rect 519 -575 522 -564
rect 531 -572 571 -569
rect 643 -573 646 -555
rect 460 -578 522 -575
rect 439 -636 506 -633
rect 357 -651 361 -648
rect 349 -660 353 -657
rect 358 -659 361 -651
rect 503 -656 506 -636
rect 653 -640 656 -541
rect 919 -544 987 -540
rect 671 -556 810 -552
rect 673 -569 690 -565
rect 1011 -572 1014 -534
rect 1172 -555 1175 -548
rect 1172 -558 1271 -555
rect 1172 -564 1175 -558
rect 1144 -567 1175 -564
rect 1144 -578 1147 -567
rect 1156 -575 1196 -572
rect 1268 -576 1271 -558
rect 1085 -581 1147 -578
rect 631 -643 656 -640
rect 225 -669 324 -666
rect 225 -675 228 -669
rect 197 -678 228 -675
rect 197 -689 200 -678
rect 209 -686 249 -683
rect 321 -687 324 -669
rect 138 -692 200 -689
rect 334 -689 337 -668
rect 350 -670 353 -660
rect 631 -670 634 -643
rect 350 -672 358 -670
rect 350 -673 354 -672
rect 485 -678 492 -675
rect 485 -684 488 -678
rect 453 -687 488 -684
rect 492 -693 497 -692
rect 453 -696 497 -693
rect 620 -687 623 -686
rect 588 -690 623 -687
rect 18 -704 41 -700
rect 22 -775 26 -704
rect 453 -705 501 -702
rect 597 -700 622 -697
rect 335 -717 338 -715
rect 307 -720 338 -717
rect 335 -726 338 -720
rect 510 -719 513 -715
rect 639 -717 642 -707
rect 663 -717 666 -625
rect 677 -641 680 -614
rect 815 -630 818 -599
rect 974 -630 977 -594
rect 815 -633 977 -630
rect 677 -644 731 -641
rect 728 -685 731 -644
rect 815 -717 818 -633
rect 829 -701 833 -672
rect 639 -719 818 -717
rect 510 -720 818 -719
rect 510 -722 642 -720
rect 510 -726 513 -722
rect 335 -729 513 -726
<< labels >>
rlabel metal1 40 55 45 58 4 VDD
rlabel metal1 40 0 45 3 2 GND
rlabel metal1 40 159 44 163 4 VDD
rlabel metal1 40 62 44 66 2 GND
rlabel metal1 -1 103 3 107 3 A0
rlabel metal1 -1 95 3 99 3 B0
rlabel metal1 144 19 148 23 1 G0
rlabel metal1 333 115 337 119 7 P0
rlabel metal1 349 116 354 119 4 VDD
rlabel metal1 349 61 354 64 2 GND
rlabel metal1 -1 178 4 183 4 Cin
rlabel metal1 467 116 470 119 4 VDD
rlabel metal1 467 61 470 64 2 GND
rlabel metal1 581 80 585 84 7 C1
rlabel metal1 291 247 295 251 4 VDD
rlabel metal1 291 150 295 154 2 GND
rlabel metal1 584 203 588 207 7 S0
rlabel metal1 39 -125 44 -122 4 VDD
rlabel metal1 39 -180 44 -177 2 GND
rlabel metal1 39 -21 43 -17 4 VDD
rlabel metal1 39 -118 43 -114 2 GND
rlabel metal1 -2 -77 2 -73 3 A1
rlabel metal1 -2 -85 2 -81 3 B1
rlabel metal1 143 -161 147 -157 1 G1
rlabel metal1 332 -65 336 -61 1 P1
rlabel metal1 355 -63 358 -60 4 VDD
rlabel metal1 355 -118 358 -115 2 GND
rlabel metal1 272 30 277 33 4 VDD
rlabel metal1 272 -25 277 -22 2 GND
rlabel metal1 396 23 399 26 4 VDD
rlabel metal1 424 -32 427 -29 1 GND
rlabel metal1 529 -13 533 -9 1 C2
rlabel metal1 171 -148 175 -144 4 VDD
rlabel metal1 171 -245 175 -241 2 GND
rlabel metal1 39 -379 44 -376 4 VDD
rlabel metal1 39 -434 44 -431 2 GND
rlabel metal1 39 -275 43 -271 4 VDD
rlabel metal1 39 -372 43 -368 2 GND
rlabel metal1 360 -301 363 -298 4 VDD
rlabel metal1 360 -356 363 -353 2 GND
rlabel metal1 -2 -331 2 -327 3 A2
rlabel metal1 -2 -339 2 -335 3 B2
rlabel metal1 329 -319 333 -315 1 P2
rlabel metal1 143 -415 147 -411 1 G2
rlabel metal1 529 -300 532 -297 4 VDD
rlabel metal1 529 -355 532 -352 2 GND
rlabel metal1 540 -280 543 -260 3 VDD
rlabel metal1 529 -236 534 -233 4 VDD
rlabel metal1 529 -291 534 -288 2 GND
rlabel metal1 676 -288 679 -285 4 VDD
rlabel metal1 676 -344 679 -341 2 GND
rlabel metal1 830 -325 834 -321 7 C3
rlabel metal1 530 -205 534 -201 2 GND
rlabel metal1 530 -108 534 -104 4 VDD
rlabel metal1 40 -561 45 -558 4 VDD
rlabel metal1 40 -616 45 -613 2 GND
rlabel metal1 40 -457 44 -453 4 VDD
rlabel metal1 40 -554 44 -550 2 GND
rlabel metal1 288 -477 291 -474 2 GND
rlabel metal1 144 -597 148 -593 1 G3
rlabel metal1 299 -413 304 -410 1 VDD
rlabel metal1 424 -412 427 -409 4 VDD
rlabel metal1 439 -467 454 -464 1 GND
rlabel metal1 570 -412 573 -409 4 VDD
rlabel metal1 597 -467 602 -464 1 GND
rlabel metal1 717 -401 720 -381 3 VDD
rlabel metal1 706 -357 711 -354 4 VDD
rlabel metal1 706 -412 711 -409 2 GND
rlabel metal1 716 -433 719 -430 4 VDD
rlabel metal1 739 -502 747 -499 1 GND
rlabel metal1 363 -526 367 -522 4 VDD
rlabel metal1 363 -623 367 -619 2 GND
rlabel metal1 333 -501 337 -497 1 P3
rlabel metal1 -1 -513 3 -509 3 A3
rlabel metal1 -1 -521 3 -517 3 B3
rlabel metal1 41 -744 46 -741 4 VDD
rlabel metal1 41 -799 46 -796 2 GND
rlabel metal1 41 -640 45 -636 4 VDD
rlabel metal1 41 -737 45 -733 2 GND
rlabel metal1 0 -696 4 -692 3 A4
rlabel metal1 0 -704 4 -700 3 B4
rlabel metal1 145 -780 149 -776 1 G4
rlabel metal1 380 -722 384 -718 1 VDD
rlabel metal1 468 -715 472 -711 1 GND
rlabel metal1 288 -708 292 -704 1 P4
rlabel metal1 506 -651 509 -648 4 VDD
rlabel metal1 532 -715 558 -712 1 GND
rlabel metal1 634 -715 637 -712 2 GND
rlabel metal1 634 -660 637 -657 4 VDD
rlabel metal1 687 -580 690 -577 4 VDD
rlabel metal1 710 -635 733 -632 1 GND
rlabel metal1 844 -601 847 -581 3 VDD
rlabel metal1 833 -557 838 -554 4 VDD
rlabel metal1 833 -612 838 -609 2 GND
rlabel metal1 1032 -717 1036 -713 1 GND
rlabel metal1 854 -718 858 -714 1 VDD
rlabel metal1 988 -529 992 -525 4 VDD
rlabel metal1 988 -626 992 -622 2 GND
rlabel metal1 1281 -573 1285 -569 7 S4
rlabel metal1 888 -469 892 -465 7 C4
rlabel metal1 1281 -509 1285 -505 7 S3
rlabel metal1 1281 -500 1285 -496 7 S2
rlabel metal1 1281 -489 1285 -485 7 S1
rlabel metal1 1280 -469 1284 -465 7 S0
rlabel metal1 1282 -582 1286 -578 7 Cout
<< end >>
