* NGSPICE file created from NAND4.ext - technology: scmos

.global Vdd Gnd 


* Top level circuit NAND4

M1000 VDD D OUT w_n6_46# cmosp w=20u l=2u
+  ad=320p pd=152u as=240p ps=104u
M1001 OUT D a_23_0# Gnd cmosn w=40u l=2u
+  ad=200p pd=90u as=240p ps=92u
M1002 OUT A VDD w_n6_46# cmosp w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_15_0# B a_7_0# Gnd cmosn w=40u l=2u
+  ad=240p pd=92u as=240p ps=92u
M1004 VDD B OUT w_n6_46# cmosp w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1005 a_7_0# A GND Gnd cmosn w=40u l=2u
+  ad=0p pd=0u as=200p ps=90u
M1006 a_23_0# C a_15_0# Gnd cmosn w=40u l=2u
+  ad=0p pd=0u as=0p ps=0u
M1007 OUT C VDD w_n6_46# cmosp w=20u l=2u
+  ad=0p pd=0u as=0p ps=0u
.end

