magic
tech scmos
timestamp 1764715846
<< nwell >>
rect 63 119 95 151
rect -28 85 4 117
rect 63 63 95 95
rect 159 85 191 117
rect -43 5 -11 37
rect 30 26 54 58
<< ntransistor >>
rect 105 138 125 140
rect 105 130 125 132
rect 14 104 34 106
rect 201 104 221 106
rect 14 96 34 98
rect 201 96 221 98
rect 105 82 125 84
rect 105 74 125 76
rect -4 24 16 26
rect -4 16 16 18
rect 41 6 43 16
<< ptransistor >>
rect 69 138 89 140
rect 69 130 89 132
rect -22 104 -2 106
rect 165 104 185 106
rect -22 96 -2 98
rect 165 96 185 98
rect 69 82 89 84
rect 69 74 89 76
rect 41 32 43 52
rect -37 24 -17 26
rect -37 16 -17 18
<< ndiffusion >>
rect 105 140 125 141
rect 105 137 125 138
rect 105 132 125 133
rect 105 129 125 130
rect 14 106 34 107
rect 14 103 34 104
rect 201 106 221 107
rect 14 98 34 99
rect 14 95 34 96
rect 201 103 221 104
rect 201 98 221 99
rect 201 95 221 96
rect 105 84 125 85
rect 105 81 125 82
rect 105 76 125 77
rect 105 73 125 74
rect -4 26 16 27
rect -4 23 16 24
rect -4 18 16 19
rect -4 15 16 16
rect 40 6 41 16
rect 43 6 44 16
<< pdiffusion >>
rect 69 140 89 141
rect 69 137 89 138
rect 69 132 89 133
rect 69 129 89 130
rect -22 106 -2 107
rect -22 103 -2 104
rect -22 98 -2 99
rect 165 106 185 107
rect 165 103 185 104
rect -22 95 -2 96
rect 165 98 185 99
rect 165 95 185 96
rect 69 84 89 85
rect 69 81 89 82
rect 69 76 89 77
rect 69 73 89 74
rect 40 32 41 52
rect 43 32 44 52
rect -37 26 -17 27
rect -37 23 -17 24
rect -37 18 -17 19
rect -37 15 -17 16
<< ndcontact >>
rect 105 141 125 145
rect 105 133 125 137
rect 105 125 125 129
rect 14 107 34 111
rect 201 107 221 111
rect 14 99 34 103
rect 201 99 221 103
rect 14 91 34 95
rect 201 91 221 95
rect 105 85 125 89
rect 105 77 125 81
rect 105 69 125 73
rect -4 27 16 31
rect -4 19 16 23
rect -4 11 16 15
rect 36 6 40 16
rect 44 6 48 16
<< pdcontact >>
rect 69 141 89 145
rect 69 133 89 137
rect 69 125 89 129
rect -22 107 -2 111
rect 165 107 185 111
rect -22 99 -2 103
rect 165 99 185 103
rect -22 91 -2 95
rect 165 91 185 95
rect 69 85 89 89
rect 69 77 89 81
rect 69 69 89 73
rect 36 32 40 52
rect 44 32 48 52
rect -37 27 -17 31
rect -37 19 -17 23
rect -37 11 -17 15
<< polysilicon >>
rect 57 138 69 140
rect 89 138 105 140
rect 125 138 128 140
rect 57 130 69 132
rect 89 130 105 132
rect 125 130 128 132
rect -34 104 -22 106
rect -2 104 14 106
rect 34 104 37 106
rect 153 104 165 106
rect 185 104 201 106
rect 221 104 224 106
rect -34 96 -22 98
rect -2 96 14 98
rect 34 96 37 98
rect 153 96 165 98
rect 185 96 201 98
rect 221 96 224 98
rect 57 82 69 84
rect 89 82 105 84
rect 125 82 128 84
rect 57 74 69 76
rect 89 74 105 76
rect 125 74 128 76
rect 41 52 43 55
rect -46 24 -37 26
rect -17 24 -4 26
rect 16 24 19 26
rect -46 16 -37 18
rect -17 16 -4 18
rect 16 16 19 18
rect 41 16 43 32
rect 41 3 43 6
<< polycontact >>
rect 53 137 57 141
rect 53 129 57 133
rect -38 103 -34 107
rect -38 95 -34 99
rect 149 103 153 107
rect 149 95 153 99
rect 53 81 57 85
rect 53 73 57 77
rect -50 23 -46 27
rect -50 15 -46 19
rect 37 19 41 23
<< metal1 >>
rect -54 159 159 163
rect 97 148 140 152
rect 60 141 69 145
rect -42 137 53 141
rect -42 107 -38 137
rect 49 118 53 133
rect 60 129 63 141
rect 97 137 101 148
rect 125 141 128 145
rect 89 133 101 137
rect 97 129 101 133
rect 6 114 53 118
rect -31 107 -22 111
rect -95 103 -38 107
rect -95 95 -82 99
rect -65 27 -61 103
rect -49 95 -38 99
rect -31 95 -28 107
rect 6 103 10 114
rect 34 107 38 111
rect -2 99 10 103
rect 6 95 10 99
rect -42 77 -38 95
rect -31 91 -22 95
rect 6 91 14 95
rect 49 81 53 114
rect 60 125 69 129
rect 97 125 105 129
rect 60 116 64 125
rect 60 112 109 116
rect 60 89 64 112
rect 136 107 140 148
rect 155 116 159 159
rect 193 115 243 119
rect 156 107 165 111
rect 136 103 149 107
rect 136 96 149 99
rect 97 95 149 96
rect 156 95 159 107
rect 193 103 197 115
rect 221 107 225 111
rect 185 99 197 103
rect 193 95 197 99
rect 97 92 140 95
rect 60 85 69 89
rect -42 73 53 77
rect 60 73 63 85
rect 97 81 101 92
rect 156 91 165 95
rect 193 91 201 95
rect 125 85 135 89
rect 89 77 101 81
rect 97 73 101 77
rect 60 69 69 73
rect 97 69 105 73
rect 131 66 135 85
rect 225 66 229 107
rect -54 62 229 66
rect -54 55 40 58
rect -43 31 -40 55
rect 36 52 40 55
rect -11 34 29 38
rect -11 31 -7 34
rect -43 27 -37 31
rect -11 27 -4 31
rect -65 23 -50 27
rect -73 15 -50 19
rect -43 15 -40 27
rect -11 23 -7 27
rect 25 23 29 34
rect 44 23 48 32
rect -17 19 -7 23
rect 25 19 37 23
rect 44 19 54 23
rect 44 16 48 19
rect -43 11 -37 15
rect 16 11 22 15
rect 19 3 22 11
rect 36 3 40 6
rect -54 0 40 3
<< m2contact >>
rect -32 154 -27 159
rect 128 140 133 145
rect -32 111 -27 116
rect -82 95 -77 100
rect -54 95 -49 100
rect 38 106 43 111
rect 109 112 114 117
rect 154 111 159 116
rect 225 107 230 112
rect -73 19 -68 24
<< metal2 >>
rect -31 116 -28 154
rect 130 133 133 140
rect 130 130 229 133
rect 130 124 133 130
rect 102 121 133 124
rect 102 110 105 121
rect 114 113 154 116
rect 226 112 229 130
rect 43 107 105 110
rect -77 95 -54 99
rect -73 24 -69 95
<< labels >>
rlabel metal1 -54 55 -49 58 4 VDD
rlabel metal1 -54 0 -49 3 2 GND
rlabel metal1 -54 159 -50 163 4 VDD
rlabel metal1 -54 62 -50 66 2 GND
rlabel metal1 -95 95 -91 99 3 B
rlabel metal1 -95 103 -91 107 3 A
rlabel metal1 50 19 54 23 1 G
rlabel metal1 239 115 243 119 7 P
<< end >>
