module AND6(input A, input B, input C, input D, input E, input F, output Y);
    assign Y = A & B & C & D & E & F;
endmodule
