magic
tech scmos
timestamp 1763742894
<< nwell >>
rect 2 -12 34 28
<< ntransistor >>
rect 40 15 70 17
rect 40 7 70 9
rect 40 -1 70 1
<< ptransistor >>
rect 8 15 28 17
rect 8 7 28 9
rect 8 -1 28 1
<< ndiffusion >>
rect 40 17 70 18
rect 40 14 70 15
rect 40 9 70 10
rect 40 6 70 7
rect 40 1 70 2
rect 40 -2 70 -1
<< pdiffusion >>
rect 8 17 28 18
rect 8 14 28 15
rect 8 9 28 10
rect 8 6 28 7
rect 8 1 28 2
rect 8 -2 28 -1
<< ndcontact >>
rect 40 18 70 22
rect 40 10 70 14
rect 40 2 70 6
rect 40 -6 70 -2
<< pdcontact >>
rect 8 18 28 22
rect 8 10 28 14
rect 8 2 28 6
rect 8 -6 28 -2
<< polysilicon >>
rect -1 15 8 17
rect 28 15 40 17
rect 70 15 73 17
rect -1 7 8 9
rect 28 7 40 9
rect 70 7 73 9
rect -1 -1 8 1
rect 28 -1 40 1
rect 70 -1 73 1
<< polycontact >>
rect -5 14 -1 18
rect -5 6 -1 10
rect -5 -2 -1 2
<< metal1 >>
rect -9 14 -5 18
rect 2 14 5 28
rect 34 25 79 28
rect 34 22 37 25
rect 28 18 40 22
rect 2 10 8 14
rect -9 6 -5 10
rect -9 -2 -5 2
rect 2 -2 5 10
rect 33 6 37 18
rect 28 2 37 6
rect 73 -2 76 22
rect 2 -6 8 -2
rect 70 -6 76 -2
rect 2 -12 5 -6
<< labels >>
rlabel metal1 73 -6 76 22 7 GND
rlabel metal1 2 -12 5 28 3 VDD
rlabel metal1 -9 -2 -5 2 3 A
rlabel metal1 -9 6 -5 10 3 B
rlabel metal1 -9 14 -5 18 3 C
rlabel metal1 76 25 79 28 6 OUT
<< end >>
