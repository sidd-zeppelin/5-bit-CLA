magic
tech scmos
timestamp 1763754879
<< nwell >>
rect -1587 1490 -1555 1522
rect -1481 1508 -1449 1540
rect -1260 1490 -1228 1522
rect -1154 1508 -1122 1540
rect -1683 1458 -1659 1490
rect -1632 1458 -1608 1490
rect -1587 1443 -1555 1475
rect -1481 1443 -1449 1475
rect -1355 1458 -1331 1490
rect -1305 1458 -1281 1490
rect -1260 1443 -1228 1475
rect -1154 1443 -1122 1475
rect -483 1461 -451 1493
rect -410 1482 -386 1514
rect -345 1425 -293 1457
rect -262 1447 -238 1479
rect -1587 1312 -1555 1344
rect -1481 1330 -1449 1362
rect -1260 1312 -1228 1344
rect -1154 1330 -1122 1362
rect -893 1359 -861 1391
rect -799 1367 -775 1399
rect -63 1344 -31 1376
rect -1683 1280 -1659 1312
rect -1632 1280 -1608 1312
rect -1587 1265 -1555 1297
rect -1481 1265 -1449 1297
rect -1355 1280 -1331 1312
rect -1305 1280 -1281 1312
rect -1260 1265 -1228 1297
rect -1154 1265 -1122 1297
rect -790 1283 -758 1315
rect -154 1310 -122 1342
rect -63 1288 -31 1320
rect 33 1310 65 1342
rect -881 1249 -849 1281
rect -790 1227 -758 1259
rect -694 1249 -662 1281
rect -1588 1137 -1556 1169
rect -1482 1155 -1450 1187
rect -1261 1137 -1229 1169
rect -1155 1155 -1123 1187
rect -494 1168 -462 1208
rect -412 1186 -388 1218
rect -35 1177 -3 1209
rect -1684 1105 -1660 1137
rect -1633 1105 -1609 1137
rect -1588 1090 -1556 1122
rect -1482 1090 -1450 1122
rect -1356 1105 -1332 1137
rect -1306 1105 -1282 1137
rect -1261 1090 -1229 1122
rect -1155 1090 -1123 1122
rect -487 1091 -455 1123
rect -414 1112 -390 1144
rect -126 1143 -94 1175
rect -35 1121 -3 1153
rect 61 1143 93 1175
rect -298 1054 -226 1094
rect -196 1073 -172 1105
rect -1588 962 -1556 994
rect -1482 980 -1450 1012
rect -1261 962 -1229 994
rect -1155 980 -1123 1012
rect -897 993 -865 1025
rect -803 1001 -779 1033
rect -1684 930 -1660 962
rect -1633 930 -1609 962
rect -1588 915 -1556 947
rect -1482 915 -1450 947
rect -1356 930 -1332 962
rect -1306 930 -1282 962
rect -1261 915 -1229 947
rect -1155 915 -1123 947
rect -794 917 -762 949
rect -885 883 -853 915
rect -794 861 -762 893
rect -698 883 -666 915
rect -1588 786 -1556 818
rect -1482 804 -1450 836
rect -1261 786 -1229 818
rect -1155 804 -1123 836
rect -454 810 -422 858
rect -362 833 -338 865
rect -233 809 -141 857
rect -110 830 -86 862
rect 73 858 105 890
rect -18 824 14 856
rect 73 802 105 834
rect 169 824 201 856
rect -1684 754 -1660 786
rect -1633 754 -1609 786
rect -1588 739 -1556 771
rect -1482 739 -1450 771
rect -1356 754 -1332 786
rect -1306 754 -1282 786
rect -1261 739 -1229 771
rect -1155 739 -1123 771
rect -452 745 -420 785
rect -370 763 -346 795
rect -1588 611 -1556 643
rect -1482 629 -1450 661
rect -1261 611 -1229 643
rect -1155 629 -1123 661
rect -897 635 -865 667
rect -803 643 -779 675
rect -452 667 -420 699
rect -379 688 -355 720
rect -1684 579 -1660 611
rect -1633 579 -1609 611
rect -1588 564 -1556 596
rect -1482 564 -1450 596
rect -1356 579 -1332 611
rect -1306 579 -1282 611
rect -1261 564 -1229 596
rect -1155 564 -1123 596
rect -794 559 -762 591
rect -885 525 -853 557
rect -794 503 -762 535
rect -698 525 -666 557
rect -1587 305 -1555 337
rect -1481 323 -1449 355
rect -1260 305 -1228 337
rect -1154 323 -1122 355
rect -1683 273 -1659 305
rect -1632 273 -1608 305
rect -1587 258 -1555 290
rect -1481 258 -1449 290
rect -1355 273 -1331 305
rect -1305 273 -1281 305
rect -1260 258 -1228 290
rect -1154 258 -1122 290
rect -897 188 -865 220
rect -803 196 -779 228
rect -1588 130 -1556 162
rect -1482 148 -1450 180
rect -1261 130 -1229 162
rect -1155 148 -1123 180
rect -1684 98 -1660 130
rect -1633 98 -1609 130
rect -1588 83 -1556 115
rect -1482 83 -1450 115
rect -1356 98 -1332 130
rect -1306 98 -1282 130
rect -1261 83 -1229 115
rect -1155 83 -1123 115
rect -794 112 -762 144
rect -885 78 -853 110
rect -794 56 -762 88
rect -698 78 -666 110
rect -1588 -45 -1556 -13
rect -1482 -27 -1450 5
rect -1261 -45 -1229 -13
rect -1155 -27 -1123 5
rect -1684 -77 -1660 -45
rect -1633 -77 -1609 -45
rect -1588 -92 -1556 -60
rect -1482 -92 -1450 -60
rect -1356 -77 -1332 -45
rect -1306 -77 -1282 -45
rect -1261 -92 -1229 -60
rect -1155 -92 -1123 -60
rect -1588 -221 -1556 -189
rect -1482 -203 -1450 -171
rect -1261 -221 -1229 -189
rect -1155 -203 -1123 -171
rect -1684 -253 -1660 -221
rect -1633 -253 -1609 -221
rect -1588 -268 -1556 -236
rect -1482 -268 -1450 -236
rect -1356 -253 -1332 -221
rect -1306 -253 -1282 -221
rect -1261 -268 -1229 -236
rect -1155 -268 -1123 -236
rect -897 -315 -865 -283
rect -803 -307 -779 -275
rect -1588 -396 -1556 -364
rect -1482 -378 -1450 -346
rect -1261 -396 -1229 -364
rect -1155 -378 -1123 -346
rect -794 -391 -762 -359
rect -1684 -428 -1660 -396
rect -1633 -428 -1609 -396
rect -1588 -443 -1556 -411
rect -1482 -443 -1450 -411
rect -1356 -428 -1332 -396
rect -1306 -428 -1282 -396
rect -1261 -443 -1229 -411
rect -1155 -443 -1123 -411
rect -885 -425 -853 -393
rect -794 -447 -762 -415
rect -698 -425 -666 -393
<< ntransistor >>
rect -1439 1527 -1419 1529
rect -1112 1527 -1092 1529
rect -1439 1519 -1419 1521
rect -1112 1519 -1092 1521
rect -1545 1509 -1525 1511
rect -1218 1509 -1198 1511
rect -1545 1501 -1525 1503
rect -1218 1501 -1198 1503
rect -1545 1462 -1525 1464
rect -444 1480 -424 1482
rect -444 1472 -424 1474
rect -1439 1462 -1419 1464
rect -1545 1454 -1525 1456
rect -1672 1440 -1670 1450
rect -1621 1440 -1619 1450
rect -1439 1454 -1419 1456
rect -1218 1462 -1198 1464
rect -1112 1462 -1092 1464
rect -399 1462 -397 1472
rect -1218 1454 -1198 1456
rect -1344 1440 -1342 1450
rect -1294 1440 -1292 1450
rect -1112 1454 -1092 1456
rect -287 1444 -277 1446
rect -287 1436 -277 1438
rect -251 1427 -249 1437
rect -851 1378 -831 1380
rect -851 1370 -831 1372
rect -21 1363 -1 1365
rect -1439 1349 -1419 1351
rect -1112 1349 -1092 1351
rect -788 1349 -786 1359
rect -21 1355 -1 1357
rect -1439 1341 -1419 1343
rect -1112 1341 -1092 1343
rect -1545 1331 -1525 1333
rect -1218 1331 -1198 1333
rect -1545 1323 -1525 1325
rect -112 1329 -92 1331
rect -1218 1323 -1198 1325
rect 75 1329 95 1331
rect -112 1321 -92 1323
rect 75 1321 95 1323
rect -1545 1284 -1525 1286
rect -21 1307 -1 1309
rect -748 1302 -728 1304
rect -21 1299 -1 1301
rect -748 1294 -728 1296
rect -1439 1284 -1419 1286
rect -1545 1276 -1525 1278
rect -1672 1262 -1670 1272
rect -1621 1262 -1619 1272
rect -1439 1276 -1419 1278
rect -1218 1284 -1198 1286
rect -1112 1284 -1092 1286
rect -1218 1276 -1198 1278
rect -1344 1262 -1342 1272
rect -1294 1262 -1292 1272
rect -1112 1276 -1092 1278
rect -839 1268 -819 1270
rect -652 1268 -632 1270
rect -839 1260 -819 1262
rect -652 1260 -632 1262
rect -748 1246 -728 1248
rect -748 1238 -728 1240
rect -456 1195 -426 1197
rect 7 1196 27 1198
rect -456 1187 -426 1189
rect -1440 1174 -1420 1176
rect -456 1179 -426 1181
rect -1113 1174 -1093 1176
rect 7 1188 27 1190
rect -1440 1166 -1420 1168
rect -1113 1166 -1093 1168
rect -401 1166 -399 1176
rect -1546 1156 -1526 1158
rect -84 1162 -64 1164
rect -1219 1156 -1199 1158
rect -1546 1148 -1526 1150
rect 103 1162 123 1164
rect -84 1154 -64 1156
rect -1219 1148 -1199 1150
rect 103 1154 123 1156
rect 7 1140 27 1142
rect -1546 1109 -1526 1111
rect 7 1132 27 1134
rect -1440 1109 -1420 1111
rect -1546 1101 -1526 1103
rect -1673 1087 -1671 1097
rect -1622 1087 -1620 1097
rect -1440 1101 -1420 1103
rect -1219 1109 -1199 1111
rect -1113 1109 -1093 1111
rect -448 1110 -428 1112
rect -1219 1101 -1199 1103
rect -1345 1087 -1343 1097
rect -1295 1087 -1293 1097
rect -1113 1101 -1093 1103
rect -448 1102 -428 1104
rect -403 1092 -401 1102
rect -220 1081 -210 1083
rect -220 1073 -210 1075
rect -220 1065 -210 1067
rect -185 1053 -183 1063
rect -855 1012 -835 1014
rect -1440 999 -1420 1001
rect -855 1004 -835 1006
rect -1113 999 -1093 1001
rect -1440 991 -1420 993
rect -1113 991 -1093 993
rect -1546 981 -1526 983
rect -792 983 -790 993
rect -1219 981 -1199 983
rect -1546 973 -1526 975
rect -1219 973 -1199 975
rect -1546 934 -1526 936
rect -1440 934 -1420 936
rect -1546 926 -1526 928
rect -1673 912 -1671 922
rect -1622 912 -1620 922
rect -1440 926 -1420 928
rect -1219 934 -1199 936
rect -1113 934 -1093 936
rect -752 936 -732 938
rect -1219 926 -1199 928
rect -1345 912 -1343 922
rect -1295 912 -1293 922
rect -1113 926 -1093 928
rect -752 928 -732 930
rect -843 902 -823 904
rect -656 902 -636 904
rect -843 894 -823 896
rect -656 894 -636 896
rect -752 880 -732 882
rect 115 877 135 879
rect -752 872 -732 874
rect 115 869 135 871
rect -416 845 -376 847
rect -135 844 -125 846
rect -416 837 -376 839
rect -1440 823 -1420 825
rect -416 829 -376 831
rect -1113 823 -1093 825
rect -1440 815 -1420 817
rect -135 836 -125 838
rect 24 843 44 845
rect -135 828 -125 830
rect -416 821 -376 823
rect -1113 815 -1093 817
rect -1546 805 -1526 807
rect -351 813 -349 823
rect -135 820 -125 822
rect 211 843 231 845
rect 24 835 44 837
rect 211 835 231 837
rect 115 821 135 823
rect -99 810 -97 820
rect 115 813 135 815
rect -1219 805 -1199 807
rect -1546 797 -1526 799
rect -1219 797 -1199 799
rect -1546 758 -1526 760
rect -414 772 -384 774
rect -1440 758 -1420 760
rect -1546 750 -1526 752
rect -1673 736 -1671 746
rect -1622 736 -1620 746
rect -1440 750 -1420 752
rect -1219 758 -1199 760
rect -414 764 -384 766
rect -1113 758 -1093 760
rect -1219 750 -1199 752
rect -1345 736 -1343 746
rect -1295 736 -1293 746
rect -414 756 -384 758
rect -1113 750 -1093 752
rect -359 743 -357 753
rect -413 686 -393 688
rect -413 678 -393 680
rect -1440 648 -1420 650
rect -855 654 -835 656
rect -1113 648 -1093 650
rect -1440 640 -1420 642
rect -368 668 -366 678
rect -855 646 -835 648
rect -1113 640 -1093 642
rect -1546 630 -1526 632
rect -1219 630 -1199 632
rect -1546 622 -1526 624
rect -792 625 -790 635
rect -1219 622 -1199 624
rect -1546 583 -1526 585
rect -1440 583 -1420 585
rect -1546 575 -1526 577
rect -1673 561 -1671 571
rect -1622 561 -1620 571
rect -1440 575 -1420 577
rect -1219 583 -1199 585
rect -1113 583 -1093 585
rect -1219 575 -1199 577
rect -1345 561 -1343 571
rect -1295 561 -1293 571
rect -752 578 -732 580
rect -1113 575 -1093 577
rect -752 570 -732 572
rect -843 544 -823 546
rect -656 544 -636 546
rect -843 536 -823 538
rect -656 536 -636 538
rect -752 522 -732 524
rect -752 514 -732 516
rect -1439 342 -1419 344
rect -1112 342 -1092 344
rect -1439 334 -1419 336
rect -1112 334 -1092 336
rect -1545 324 -1525 326
rect -1218 324 -1198 326
rect -1545 316 -1525 318
rect -1218 316 -1198 318
rect -1545 277 -1525 279
rect -1439 277 -1419 279
rect -1545 269 -1525 271
rect -1672 255 -1670 265
rect -1621 255 -1619 265
rect -1439 269 -1419 271
rect -1218 277 -1198 279
rect -1112 277 -1092 279
rect -1218 269 -1198 271
rect -1344 255 -1342 265
rect -1294 255 -1292 265
rect -1112 269 -1092 271
rect -855 207 -835 209
rect -855 199 -835 201
rect -792 178 -790 188
rect -1440 167 -1420 169
rect -1113 167 -1093 169
rect -1440 159 -1420 161
rect -1113 159 -1093 161
rect -1546 149 -1526 151
rect -1219 149 -1199 151
rect -1546 141 -1526 143
rect -1219 141 -1199 143
rect -752 131 -732 133
rect -1546 102 -1526 104
rect -752 123 -732 125
rect -1440 102 -1420 104
rect -1546 94 -1526 96
rect -1673 80 -1671 90
rect -1622 80 -1620 90
rect -1440 94 -1420 96
rect -1219 102 -1199 104
rect -1113 102 -1093 104
rect -1219 94 -1199 96
rect -1345 80 -1343 90
rect -1295 80 -1293 90
rect -843 97 -823 99
rect -1113 94 -1093 96
rect -656 97 -636 99
rect -843 89 -823 91
rect -656 89 -636 91
rect -752 75 -732 77
rect -752 67 -732 69
rect -1440 -8 -1420 -6
rect -1113 -8 -1093 -6
rect -1440 -16 -1420 -14
rect -1113 -16 -1093 -14
rect -1546 -26 -1526 -24
rect -1219 -26 -1199 -24
rect -1546 -34 -1526 -32
rect -1219 -34 -1199 -32
rect -1546 -73 -1526 -71
rect -1440 -73 -1420 -71
rect -1546 -81 -1526 -79
rect -1673 -95 -1671 -85
rect -1622 -95 -1620 -85
rect -1440 -81 -1420 -79
rect -1219 -73 -1199 -71
rect -1113 -73 -1093 -71
rect -1219 -81 -1199 -79
rect -1345 -95 -1343 -85
rect -1295 -95 -1293 -85
rect -1113 -81 -1093 -79
rect -1440 -184 -1420 -182
rect -1113 -184 -1093 -182
rect -1440 -192 -1420 -190
rect -1113 -192 -1093 -190
rect -1546 -202 -1526 -200
rect -1219 -202 -1199 -200
rect -1546 -210 -1526 -208
rect -1219 -210 -1199 -208
rect -1546 -249 -1526 -247
rect -1440 -249 -1420 -247
rect -1546 -257 -1526 -255
rect -1673 -271 -1671 -261
rect -1622 -271 -1620 -261
rect -1440 -257 -1420 -255
rect -1219 -249 -1199 -247
rect -1113 -249 -1093 -247
rect -1219 -257 -1199 -255
rect -1345 -271 -1343 -261
rect -1295 -271 -1293 -261
rect -1113 -257 -1093 -255
rect -855 -296 -835 -294
rect -855 -304 -835 -302
rect -792 -325 -790 -315
rect -1440 -359 -1420 -357
rect -1113 -359 -1093 -357
rect -1440 -367 -1420 -365
rect -1113 -367 -1093 -365
rect -1546 -377 -1526 -375
rect -752 -372 -732 -370
rect -1219 -377 -1199 -375
rect -1546 -385 -1526 -383
rect -752 -380 -732 -378
rect -1219 -385 -1199 -383
rect -1546 -424 -1526 -422
rect -843 -406 -823 -404
rect -656 -406 -636 -404
rect -843 -414 -823 -412
rect -1440 -424 -1420 -422
rect -1546 -432 -1526 -430
rect -1673 -446 -1671 -436
rect -1622 -446 -1620 -436
rect -1440 -432 -1420 -430
rect -1219 -424 -1199 -422
rect -656 -414 -636 -412
rect -1113 -424 -1093 -422
rect -1219 -432 -1199 -430
rect -1345 -446 -1343 -436
rect -1295 -446 -1293 -436
rect -752 -428 -732 -426
rect -1113 -432 -1093 -430
rect -752 -436 -732 -434
<< ptransistor >>
rect -1475 1527 -1455 1529
rect -1148 1527 -1128 1529
rect -1475 1519 -1455 1521
rect -1148 1519 -1128 1521
rect -1581 1509 -1561 1511
rect -1254 1509 -1234 1511
rect -1581 1501 -1561 1503
rect -1254 1501 -1234 1503
rect -399 1488 -397 1508
rect -1672 1464 -1670 1484
rect -1621 1464 -1619 1484
rect -1581 1462 -1561 1464
rect -1344 1464 -1342 1484
rect -1294 1464 -1292 1484
rect -477 1480 -457 1482
rect -477 1472 -457 1474
rect -1475 1462 -1455 1464
rect -1581 1454 -1561 1456
rect -1475 1454 -1455 1456
rect -1254 1462 -1234 1464
rect -1148 1462 -1128 1464
rect -1254 1454 -1234 1456
rect -1148 1454 -1128 1456
rect -251 1453 -249 1473
rect -339 1444 -299 1446
rect -339 1436 -299 1438
rect -887 1378 -867 1380
rect -788 1373 -786 1393
rect -887 1370 -867 1372
rect -57 1363 -37 1365
rect -1475 1349 -1455 1351
rect -1148 1349 -1128 1351
rect -57 1355 -37 1357
rect -1475 1341 -1455 1343
rect -1148 1341 -1128 1343
rect -1581 1331 -1561 1333
rect -1254 1331 -1234 1333
rect -1581 1323 -1561 1325
rect -148 1329 -128 1331
rect -1254 1323 -1234 1325
rect 39 1329 59 1331
rect -148 1321 -128 1323
rect 39 1321 59 1323
rect -1672 1286 -1670 1306
rect -1621 1286 -1619 1306
rect -1581 1284 -1561 1286
rect -1344 1286 -1342 1306
rect -1294 1286 -1292 1306
rect -57 1307 -37 1309
rect -784 1302 -764 1304
rect -57 1299 -37 1301
rect -784 1294 -764 1296
rect -1475 1284 -1455 1286
rect -1581 1276 -1561 1278
rect -1475 1276 -1455 1278
rect -1254 1284 -1234 1286
rect -1148 1284 -1128 1286
rect -1254 1276 -1234 1278
rect -1148 1276 -1128 1278
rect -875 1268 -855 1270
rect -688 1268 -668 1270
rect -875 1260 -855 1262
rect -688 1260 -668 1262
rect -784 1246 -764 1248
rect -784 1238 -764 1240
rect -488 1195 -468 1197
rect -401 1192 -399 1212
rect -29 1196 -9 1198
rect -488 1187 -468 1189
rect -1476 1174 -1456 1176
rect -488 1179 -468 1181
rect -1149 1174 -1129 1176
rect -29 1188 -9 1190
rect -1476 1166 -1456 1168
rect -1149 1166 -1129 1168
rect -1582 1156 -1562 1158
rect -120 1162 -100 1164
rect -1255 1156 -1235 1158
rect -1582 1148 -1562 1150
rect 67 1162 87 1164
rect -120 1154 -100 1156
rect -1255 1148 -1235 1150
rect 67 1154 87 1156
rect -29 1140 -9 1142
rect -1673 1111 -1671 1131
rect -1622 1111 -1620 1131
rect -1582 1109 -1562 1111
rect -1345 1111 -1343 1131
rect -1295 1111 -1293 1131
rect -403 1118 -401 1138
rect -29 1132 -9 1134
rect -1476 1109 -1456 1111
rect -1582 1101 -1562 1103
rect -1476 1101 -1456 1103
rect -1255 1109 -1235 1111
rect -1149 1109 -1129 1111
rect -481 1110 -461 1112
rect -1255 1101 -1235 1103
rect -1149 1101 -1129 1103
rect -481 1102 -461 1104
rect -292 1081 -232 1083
rect -185 1079 -183 1099
rect -292 1073 -232 1075
rect -292 1065 -232 1067
rect -891 1012 -871 1014
rect -1476 999 -1456 1001
rect -792 1007 -790 1027
rect -891 1004 -871 1006
rect -1149 999 -1129 1001
rect -1476 991 -1456 993
rect -1149 991 -1129 993
rect -1582 981 -1562 983
rect -1255 981 -1235 983
rect -1582 973 -1562 975
rect -1255 973 -1235 975
rect -1673 936 -1671 956
rect -1622 936 -1620 956
rect -1582 934 -1562 936
rect -1345 936 -1343 956
rect -1295 936 -1293 956
rect -1476 934 -1456 936
rect -1582 926 -1562 928
rect -1476 926 -1456 928
rect -1255 934 -1235 936
rect -1149 934 -1129 936
rect -788 936 -768 938
rect -1255 926 -1235 928
rect -1149 926 -1129 928
rect -788 928 -768 930
rect -879 902 -859 904
rect -692 902 -672 904
rect -879 894 -859 896
rect -692 894 -672 896
rect -788 880 -768 882
rect 79 877 99 879
rect -788 872 -768 874
rect 79 869 99 871
rect -448 845 -428 847
rect -351 839 -349 859
rect -227 844 -147 846
rect -448 837 -428 839
rect -1476 823 -1456 825
rect -448 829 -428 831
rect -1149 823 -1129 825
rect -1476 815 -1456 817
rect -227 836 -147 838
rect -99 836 -97 856
rect -12 843 8 845
rect -227 828 -147 830
rect -448 821 -428 823
rect -1149 815 -1129 817
rect -1582 805 -1562 807
rect -227 820 -147 822
rect 175 843 195 845
rect -12 835 8 837
rect 175 835 195 837
rect 79 821 99 823
rect 79 813 99 815
rect -1255 805 -1235 807
rect -1582 797 -1562 799
rect -1255 797 -1235 799
rect -1673 760 -1671 780
rect -1622 760 -1620 780
rect -1582 758 -1562 760
rect -1345 760 -1343 780
rect -1295 760 -1293 780
rect -446 772 -426 774
rect -1476 758 -1456 760
rect -1582 750 -1562 752
rect -1476 750 -1456 752
rect -1255 758 -1235 760
rect -359 769 -357 789
rect -446 764 -426 766
rect -1149 758 -1129 760
rect -1255 750 -1235 752
rect -446 756 -426 758
rect -1149 750 -1129 752
rect -368 694 -366 714
rect -446 686 -426 688
rect -446 678 -426 680
rect -1476 648 -1456 650
rect -891 654 -871 656
rect -1149 648 -1129 650
rect -1476 640 -1456 642
rect -792 649 -790 669
rect -891 646 -871 648
rect -1149 640 -1129 642
rect -1582 630 -1562 632
rect -1255 630 -1235 632
rect -1582 622 -1562 624
rect -1255 622 -1235 624
rect -1673 585 -1671 605
rect -1622 585 -1620 605
rect -1582 583 -1562 585
rect -1345 585 -1343 605
rect -1295 585 -1293 605
rect -1476 583 -1456 585
rect -1582 575 -1562 577
rect -1476 575 -1456 577
rect -1255 583 -1235 585
rect -1149 583 -1129 585
rect -1255 575 -1235 577
rect -788 578 -768 580
rect -1149 575 -1129 577
rect -788 570 -768 572
rect -879 544 -859 546
rect -692 544 -672 546
rect -879 536 -859 538
rect -692 536 -672 538
rect -788 522 -768 524
rect -788 514 -768 516
rect -1475 342 -1455 344
rect -1148 342 -1128 344
rect -1475 334 -1455 336
rect -1148 334 -1128 336
rect -1581 324 -1561 326
rect -1254 324 -1234 326
rect -1581 316 -1561 318
rect -1254 316 -1234 318
rect -1672 279 -1670 299
rect -1621 279 -1619 299
rect -1581 277 -1561 279
rect -1344 279 -1342 299
rect -1294 279 -1292 299
rect -1475 277 -1455 279
rect -1581 269 -1561 271
rect -1475 269 -1455 271
rect -1254 277 -1234 279
rect -1148 277 -1128 279
rect -1254 269 -1234 271
rect -1148 269 -1128 271
rect -891 207 -871 209
rect -792 202 -790 222
rect -891 199 -871 201
rect -1476 167 -1456 169
rect -1149 167 -1129 169
rect -1476 159 -1456 161
rect -1149 159 -1129 161
rect -1582 149 -1562 151
rect -1255 149 -1235 151
rect -1582 141 -1562 143
rect -1255 141 -1235 143
rect -788 131 -768 133
rect -1673 104 -1671 124
rect -1622 104 -1620 124
rect -1582 102 -1562 104
rect -1345 104 -1343 124
rect -1295 104 -1293 124
rect -788 123 -768 125
rect -1476 102 -1456 104
rect -1582 94 -1562 96
rect -1476 94 -1456 96
rect -1255 102 -1235 104
rect -1149 102 -1129 104
rect -1255 94 -1235 96
rect -879 97 -859 99
rect -1149 94 -1129 96
rect -692 97 -672 99
rect -879 89 -859 91
rect -692 89 -672 91
rect -788 75 -768 77
rect -788 67 -768 69
rect -1476 -8 -1456 -6
rect -1149 -8 -1129 -6
rect -1476 -16 -1456 -14
rect -1149 -16 -1129 -14
rect -1582 -26 -1562 -24
rect -1255 -26 -1235 -24
rect -1582 -34 -1562 -32
rect -1255 -34 -1235 -32
rect -1673 -71 -1671 -51
rect -1622 -71 -1620 -51
rect -1582 -73 -1562 -71
rect -1345 -71 -1343 -51
rect -1295 -71 -1293 -51
rect -1476 -73 -1456 -71
rect -1582 -81 -1562 -79
rect -1476 -81 -1456 -79
rect -1255 -73 -1235 -71
rect -1149 -73 -1129 -71
rect -1255 -81 -1235 -79
rect -1149 -81 -1129 -79
rect -1476 -184 -1456 -182
rect -1149 -184 -1129 -182
rect -1476 -192 -1456 -190
rect -1149 -192 -1129 -190
rect -1582 -202 -1562 -200
rect -1255 -202 -1235 -200
rect -1582 -210 -1562 -208
rect -1255 -210 -1235 -208
rect -1673 -247 -1671 -227
rect -1622 -247 -1620 -227
rect -1582 -249 -1562 -247
rect -1345 -247 -1343 -227
rect -1295 -247 -1293 -227
rect -1476 -249 -1456 -247
rect -1582 -257 -1562 -255
rect -1476 -257 -1456 -255
rect -1255 -249 -1235 -247
rect -1149 -249 -1129 -247
rect -1255 -257 -1235 -255
rect -1149 -257 -1129 -255
rect -891 -296 -871 -294
rect -792 -301 -790 -281
rect -891 -304 -871 -302
rect -1476 -359 -1456 -357
rect -1149 -359 -1129 -357
rect -1476 -367 -1456 -365
rect -1149 -367 -1129 -365
rect -1582 -377 -1562 -375
rect -788 -372 -768 -370
rect -1255 -377 -1235 -375
rect -1582 -385 -1562 -383
rect -788 -380 -768 -378
rect -1255 -385 -1235 -383
rect -1673 -422 -1671 -402
rect -1622 -422 -1620 -402
rect -1582 -424 -1562 -422
rect -1345 -422 -1343 -402
rect -1295 -422 -1293 -402
rect -879 -406 -859 -404
rect -692 -406 -672 -404
rect -879 -414 -859 -412
rect -1476 -424 -1456 -422
rect -1582 -432 -1562 -430
rect -1476 -432 -1456 -430
rect -1255 -424 -1235 -422
rect -692 -414 -672 -412
rect -1149 -424 -1129 -422
rect -1255 -432 -1235 -430
rect -788 -428 -768 -426
rect -1149 -432 -1129 -430
rect -788 -436 -768 -434
<< ndiffusion >>
rect -1439 1529 -1419 1530
rect -1439 1526 -1419 1527
rect -1112 1529 -1092 1530
rect -1439 1521 -1419 1522
rect -1439 1518 -1419 1519
rect -1112 1526 -1092 1527
rect -1112 1521 -1092 1522
rect -1545 1511 -1525 1512
rect -1545 1508 -1525 1509
rect -1112 1518 -1092 1519
rect -1218 1511 -1198 1512
rect -1545 1503 -1525 1504
rect -1545 1500 -1525 1501
rect -1218 1508 -1198 1509
rect -1218 1503 -1198 1504
rect -1218 1500 -1198 1501
rect -1545 1464 -1525 1465
rect -1545 1461 -1525 1462
rect -1439 1464 -1419 1465
rect -444 1482 -424 1483
rect -444 1479 -424 1480
rect -444 1474 -424 1475
rect -1545 1456 -1525 1457
rect -1673 1440 -1672 1450
rect -1670 1440 -1669 1450
rect -1622 1440 -1621 1450
rect -1619 1440 -1618 1450
rect -1545 1453 -1525 1454
rect -1439 1461 -1419 1462
rect -1439 1456 -1419 1457
rect -1439 1453 -1419 1454
rect -1218 1464 -1198 1465
rect -1218 1461 -1198 1462
rect -444 1471 -424 1472
rect -1112 1464 -1092 1465
rect -400 1462 -399 1472
rect -397 1462 -396 1472
rect -1218 1456 -1198 1457
rect -1345 1440 -1344 1450
rect -1342 1440 -1341 1450
rect -1295 1440 -1294 1450
rect -1292 1440 -1291 1450
rect -1218 1453 -1198 1454
rect -1112 1461 -1092 1462
rect -1112 1456 -1092 1457
rect -1112 1453 -1092 1454
rect -287 1446 -277 1447
rect -287 1443 -277 1444
rect -287 1438 -277 1439
rect -287 1435 -277 1436
rect -252 1427 -251 1437
rect -249 1427 -248 1437
rect -851 1380 -831 1381
rect -851 1377 -831 1378
rect -851 1372 -831 1373
rect -851 1369 -831 1370
rect -21 1365 -1 1366
rect -1439 1351 -1419 1352
rect -1439 1348 -1419 1349
rect -1112 1351 -1092 1352
rect -789 1349 -788 1359
rect -786 1349 -785 1359
rect -21 1362 -1 1363
rect -21 1357 -1 1358
rect -21 1354 -1 1355
rect -1439 1343 -1419 1344
rect -1439 1340 -1419 1341
rect -1112 1348 -1092 1349
rect -1112 1343 -1092 1344
rect -1545 1333 -1525 1334
rect -1545 1330 -1525 1331
rect -1112 1340 -1092 1341
rect -1218 1333 -1198 1334
rect -1545 1325 -1525 1326
rect -1545 1322 -1525 1323
rect -1218 1330 -1198 1331
rect -112 1331 -92 1332
rect -1218 1325 -1198 1326
rect -1218 1322 -1198 1323
rect -112 1328 -92 1329
rect 75 1331 95 1332
rect -112 1323 -92 1324
rect -112 1320 -92 1321
rect 75 1328 95 1329
rect 75 1323 95 1324
rect 75 1320 95 1321
rect -1545 1286 -1525 1287
rect -1545 1283 -1525 1284
rect -1439 1286 -1419 1287
rect -21 1309 -1 1310
rect -748 1304 -728 1305
rect -748 1301 -728 1302
rect -21 1306 -1 1307
rect -21 1301 -1 1302
rect -748 1296 -728 1297
rect -21 1298 -1 1299
rect -1545 1278 -1525 1279
rect -1673 1262 -1672 1272
rect -1670 1262 -1669 1272
rect -1622 1262 -1621 1272
rect -1619 1262 -1618 1272
rect -1545 1275 -1525 1276
rect -1439 1283 -1419 1284
rect -1439 1278 -1419 1279
rect -1439 1275 -1419 1276
rect -1218 1286 -1198 1287
rect -1218 1283 -1198 1284
rect -748 1293 -728 1294
rect -1112 1286 -1092 1287
rect -1218 1278 -1198 1279
rect -1345 1262 -1344 1272
rect -1342 1262 -1341 1272
rect -1295 1262 -1294 1272
rect -1292 1262 -1291 1272
rect -1218 1275 -1198 1276
rect -1112 1283 -1092 1284
rect -1112 1278 -1092 1279
rect -1112 1275 -1092 1276
rect -839 1270 -819 1271
rect -839 1267 -819 1268
rect -652 1270 -632 1271
rect -839 1262 -819 1263
rect -839 1259 -819 1260
rect -652 1267 -632 1268
rect -652 1262 -632 1263
rect -652 1259 -632 1260
rect -748 1248 -728 1249
rect -748 1245 -728 1246
rect -748 1240 -728 1241
rect -748 1237 -728 1238
rect -456 1197 -426 1198
rect -456 1194 -426 1195
rect 7 1198 27 1199
rect -456 1189 -426 1190
rect -1440 1176 -1420 1177
rect -1440 1173 -1420 1174
rect -456 1186 -426 1187
rect -456 1181 -426 1182
rect -1113 1176 -1093 1177
rect -456 1178 -426 1179
rect 7 1195 27 1196
rect 7 1190 27 1191
rect 7 1187 27 1188
rect -1440 1168 -1420 1169
rect -1440 1165 -1420 1166
rect -1113 1173 -1093 1174
rect -1113 1168 -1093 1169
rect -402 1166 -401 1176
rect -399 1166 -398 1176
rect -1546 1158 -1526 1159
rect -1546 1155 -1526 1156
rect -1113 1165 -1093 1166
rect -84 1164 -64 1165
rect -1219 1158 -1199 1159
rect -1546 1150 -1526 1151
rect -1546 1147 -1526 1148
rect -1219 1155 -1199 1156
rect -84 1161 -64 1162
rect 103 1164 123 1165
rect -84 1156 -64 1157
rect -1219 1150 -1199 1151
rect -84 1153 -64 1154
rect 103 1161 123 1162
rect 103 1156 123 1157
rect 103 1153 123 1154
rect -1219 1147 -1199 1148
rect 7 1142 27 1143
rect -1546 1111 -1526 1112
rect -1546 1108 -1526 1109
rect -1440 1111 -1420 1112
rect 7 1139 27 1140
rect 7 1134 27 1135
rect 7 1131 27 1132
rect -1546 1103 -1526 1104
rect -1674 1087 -1673 1097
rect -1671 1087 -1670 1097
rect -1623 1087 -1622 1097
rect -1620 1087 -1619 1097
rect -1546 1100 -1526 1101
rect -1440 1108 -1420 1109
rect -1440 1103 -1420 1104
rect -1440 1100 -1420 1101
rect -1219 1111 -1199 1112
rect -1219 1108 -1199 1109
rect -1113 1111 -1093 1112
rect -448 1112 -428 1113
rect -1219 1103 -1199 1104
rect -1346 1087 -1345 1097
rect -1343 1087 -1342 1097
rect -1296 1087 -1295 1097
rect -1293 1087 -1292 1097
rect -1219 1100 -1199 1101
rect -1113 1108 -1093 1109
rect -1113 1103 -1093 1104
rect -448 1109 -428 1110
rect -448 1104 -428 1105
rect -1113 1100 -1093 1101
rect -448 1101 -428 1102
rect -404 1092 -403 1102
rect -401 1092 -400 1102
rect -220 1083 -210 1084
rect -220 1080 -210 1081
rect -220 1075 -210 1076
rect -220 1072 -210 1073
rect -220 1067 -210 1068
rect -220 1064 -210 1065
rect -186 1053 -185 1063
rect -183 1053 -182 1063
rect -855 1014 -835 1015
rect -1440 1001 -1420 1002
rect -1440 998 -1420 999
rect -855 1011 -835 1012
rect -855 1006 -835 1007
rect -1113 1001 -1093 1002
rect -855 1003 -835 1004
rect -1440 993 -1420 994
rect -1440 990 -1420 991
rect -1113 998 -1093 999
rect -1113 993 -1093 994
rect -1546 983 -1526 984
rect -1546 980 -1526 981
rect -1113 990 -1093 991
rect -1219 983 -1199 984
rect -793 983 -792 993
rect -790 983 -789 993
rect -1546 975 -1526 976
rect -1546 972 -1526 973
rect -1219 980 -1199 981
rect -1219 975 -1199 976
rect -1219 972 -1199 973
rect -1546 936 -1526 937
rect -1546 933 -1526 934
rect -1440 936 -1420 937
rect -1546 928 -1526 929
rect -1674 912 -1673 922
rect -1671 912 -1670 922
rect -1623 912 -1622 922
rect -1620 912 -1619 922
rect -1546 925 -1526 926
rect -1440 933 -1420 934
rect -1440 928 -1420 929
rect -1440 925 -1420 926
rect -1219 936 -1199 937
rect -1219 933 -1199 934
rect -1113 936 -1093 937
rect -752 938 -732 939
rect -1219 928 -1199 929
rect -1346 912 -1345 922
rect -1343 912 -1342 922
rect -1296 912 -1295 922
rect -1293 912 -1292 922
rect -1219 925 -1199 926
rect -1113 933 -1093 934
rect -1113 928 -1093 929
rect -752 935 -732 936
rect -752 930 -732 931
rect -1113 925 -1093 926
rect -752 927 -732 928
rect -843 904 -823 905
rect -843 901 -823 902
rect -656 904 -636 905
rect -843 896 -823 897
rect -843 893 -823 894
rect -656 901 -636 902
rect -656 896 -636 897
rect -656 893 -636 894
rect -752 882 -732 883
rect -752 879 -732 880
rect 115 879 135 880
rect -752 874 -732 875
rect -752 871 -732 872
rect 115 876 135 877
rect 115 871 135 872
rect 115 868 135 869
rect -416 847 -376 848
rect -416 844 -376 845
rect -416 839 -376 840
rect -135 846 -125 847
rect -1440 825 -1420 826
rect -1440 822 -1420 823
rect -416 836 -376 837
rect -416 831 -376 832
rect -1113 825 -1093 826
rect -1440 817 -1420 818
rect -1440 814 -1420 815
rect -1113 822 -1093 823
rect -416 828 -376 829
rect -416 823 -376 824
rect -135 843 -125 844
rect -135 838 -125 839
rect 24 845 44 846
rect -135 835 -125 836
rect -135 830 -125 831
rect -1113 817 -1093 818
rect -416 820 -376 821
rect -1546 807 -1526 808
rect -1546 804 -1526 805
rect -1113 814 -1093 815
rect -352 813 -351 823
rect -349 813 -348 823
rect -135 827 -125 828
rect -135 822 -125 823
rect 24 842 44 843
rect 211 845 231 846
rect 24 837 44 838
rect 24 834 44 835
rect 211 842 231 843
rect 211 837 231 838
rect 211 834 231 835
rect 115 823 135 824
rect -135 819 -125 820
rect -100 810 -99 820
rect -97 810 -96 820
rect 115 820 135 821
rect 115 815 135 816
rect -1219 807 -1199 808
rect 115 812 135 813
rect -1546 799 -1526 800
rect -1546 796 -1526 797
rect -1219 804 -1199 805
rect -1219 799 -1199 800
rect -1219 796 -1199 797
rect -1546 760 -1526 761
rect -1546 757 -1526 758
rect -1440 760 -1420 761
rect -414 774 -384 775
rect -1546 752 -1526 753
rect -1674 736 -1673 746
rect -1671 736 -1670 746
rect -1623 736 -1622 746
rect -1620 736 -1619 746
rect -1546 749 -1526 750
rect -1440 757 -1420 758
rect -1440 752 -1420 753
rect -1440 749 -1420 750
rect -1219 760 -1199 761
rect -1219 757 -1199 758
rect -414 771 -384 772
rect -414 766 -384 767
rect -1113 760 -1093 761
rect -1219 752 -1199 753
rect -1346 736 -1345 746
rect -1343 736 -1342 746
rect -1296 736 -1295 746
rect -1293 736 -1292 746
rect -1219 749 -1199 750
rect -1113 757 -1093 758
rect -414 763 -384 764
rect -414 758 -384 759
rect -1113 752 -1093 753
rect -414 755 -384 756
rect -1113 749 -1093 750
rect -360 743 -359 753
rect -357 743 -356 753
rect -413 688 -393 689
rect -413 685 -393 686
rect -413 680 -393 681
rect -413 677 -393 678
rect -1440 650 -1420 651
rect -1440 647 -1420 648
rect -855 656 -835 657
rect -1113 650 -1093 651
rect -1440 642 -1420 643
rect -1440 639 -1420 640
rect -1113 647 -1093 648
rect -855 653 -835 654
rect -369 668 -368 678
rect -366 668 -365 678
rect -855 648 -835 649
rect -1113 642 -1093 643
rect -855 645 -835 646
rect -1546 632 -1526 633
rect -1546 629 -1526 630
rect -1113 639 -1093 640
rect -1219 632 -1199 633
rect -1546 624 -1526 625
rect -1546 621 -1526 622
rect -1219 629 -1199 630
rect -793 625 -792 635
rect -790 625 -789 635
rect -1219 624 -1199 625
rect -1219 621 -1199 622
rect -1546 585 -1526 586
rect -1546 582 -1526 583
rect -1440 585 -1420 586
rect -1546 577 -1526 578
rect -1674 561 -1673 571
rect -1671 561 -1670 571
rect -1623 561 -1622 571
rect -1620 561 -1619 571
rect -1546 574 -1526 575
rect -1440 582 -1420 583
rect -1440 577 -1420 578
rect -1440 574 -1420 575
rect -1219 585 -1199 586
rect -1219 582 -1199 583
rect -1113 585 -1093 586
rect -1219 577 -1199 578
rect -1346 561 -1345 571
rect -1343 561 -1342 571
rect -1296 561 -1295 571
rect -1293 561 -1292 571
rect -1219 574 -1199 575
rect -1113 582 -1093 583
rect -1113 577 -1093 578
rect -752 580 -732 581
rect -1113 574 -1093 575
rect -752 577 -732 578
rect -752 572 -732 573
rect -752 569 -732 570
rect -843 546 -823 547
rect -843 543 -823 544
rect -656 546 -636 547
rect -843 538 -823 539
rect -843 535 -823 536
rect -656 543 -636 544
rect -656 538 -636 539
rect -656 535 -636 536
rect -752 524 -732 525
rect -752 521 -732 522
rect -752 516 -732 517
rect -752 513 -732 514
rect -1439 344 -1419 345
rect -1439 341 -1419 342
rect -1112 344 -1092 345
rect -1439 336 -1419 337
rect -1439 333 -1419 334
rect -1112 341 -1092 342
rect -1112 336 -1092 337
rect -1545 326 -1525 327
rect -1545 323 -1525 324
rect -1112 333 -1092 334
rect -1218 326 -1198 327
rect -1545 318 -1525 319
rect -1545 315 -1525 316
rect -1218 323 -1198 324
rect -1218 318 -1198 319
rect -1218 315 -1198 316
rect -1545 279 -1525 280
rect -1545 276 -1525 277
rect -1439 279 -1419 280
rect -1545 271 -1525 272
rect -1673 255 -1672 265
rect -1670 255 -1669 265
rect -1622 255 -1621 265
rect -1619 255 -1618 265
rect -1545 268 -1525 269
rect -1439 276 -1419 277
rect -1439 271 -1419 272
rect -1439 268 -1419 269
rect -1218 279 -1198 280
rect -1218 276 -1198 277
rect -1112 279 -1092 280
rect -1218 271 -1198 272
rect -1345 255 -1344 265
rect -1342 255 -1341 265
rect -1295 255 -1294 265
rect -1292 255 -1291 265
rect -1218 268 -1198 269
rect -1112 276 -1092 277
rect -1112 271 -1092 272
rect -1112 268 -1092 269
rect -855 209 -835 210
rect -855 206 -835 207
rect -855 201 -835 202
rect -855 198 -835 199
rect -793 178 -792 188
rect -790 178 -789 188
rect -1440 169 -1420 170
rect -1440 166 -1420 167
rect -1113 169 -1093 170
rect -1440 161 -1420 162
rect -1440 158 -1420 159
rect -1113 166 -1093 167
rect -1113 161 -1093 162
rect -1546 151 -1526 152
rect -1546 148 -1526 149
rect -1113 158 -1093 159
rect -1219 151 -1199 152
rect -1546 143 -1526 144
rect -1546 140 -1526 141
rect -1219 148 -1199 149
rect -1219 143 -1199 144
rect -1219 140 -1199 141
rect -752 133 -732 134
rect -1546 104 -1526 105
rect -1546 101 -1526 102
rect -1440 104 -1420 105
rect -752 130 -732 131
rect -752 125 -732 126
rect -752 122 -732 123
rect -1546 96 -1526 97
rect -1674 80 -1673 90
rect -1671 80 -1670 90
rect -1623 80 -1622 90
rect -1620 80 -1619 90
rect -1546 93 -1526 94
rect -1440 101 -1420 102
rect -1440 96 -1420 97
rect -1440 93 -1420 94
rect -1219 104 -1199 105
rect -1219 101 -1199 102
rect -1113 104 -1093 105
rect -1219 96 -1199 97
rect -1346 80 -1345 90
rect -1343 80 -1342 90
rect -1296 80 -1295 90
rect -1293 80 -1292 90
rect -1219 93 -1199 94
rect -1113 101 -1093 102
rect -1113 96 -1093 97
rect -843 99 -823 100
rect -1113 93 -1093 94
rect -843 96 -823 97
rect -656 99 -636 100
rect -843 91 -823 92
rect -843 88 -823 89
rect -656 96 -636 97
rect -656 91 -636 92
rect -656 88 -636 89
rect -752 77 -732 78
rect -752 74 -732 75
rect -752 69 -732 70
rect -752 66 -732 67
rect -1440 -6 -1420 -5
rect -1440 -9 -1420 -8
rect -1113 -6 -1093 -5
rect -1440 -14 -1420 -13
rect -1440 -17 -1420 -16
rect -1113 -9 -1093 -8
rect -1113 -14 -1093 -13
rect -1546 -24 -1526 -23
rect -1546 -27 -1526 -26
rect -1113 -17 -1093 -16
rect -1219 -24 -1199 -23
rect -1546 -32 -1526 -31
rect -1546 -35 -1526 -34
rect -1219 -27 -1199 -26
rect -1219 -32 -1199 -31
rect -1219 -35 -1199 -34
rect -1546 -71 -1526 -70
rect -1546 -74 -1526 -73
rect -1440 -71 -1420 -70
rect -1546 -79 -1526 -78
rect -1674 -95 -1673 -85
rect -1671 -95 -1670 -85
rect -1623 -95 -1622 -85
rect -1620 -95 -1619 -85
rect -1546 -82 -1526 -81
rect -1440 -74 -1420 -73
rect -1440 -79 -1420 -78
rect -1440 -82 -1420 -81
rect -1219 -71 -1199 -70
rect -1219 -74 -1199 -73
rect -1113 -71 -1093 -70
rect -1219 -79 -1199 -78
rect -1346 -95 -1345 -85
rect -1343 -95 -1342 -85
rect -1296 -95 -1295 -85
rect -1293 -95 -1292 -85
rect -1219 -82 -1199 -81
rect -1113 -74 -1093 -73
rect -1113 -79 -1093 -78
rect -1113 -82 -1093 -81
rect -1440 -182 -1420 -181
rect -1440 -185 -1420 -184
rect -1113 -182 -1093 -181
rect -1440 -190 -1420 -189
rect -1440 -193 -1420 -192
rect -1113 -185 -1093 -184
rect -1113 -190 -1093 -189
rect -1546 -200 -1526 -199
rect -1546 -203 -1526 -202
rect -1113 -193 -1093 -192
rect -1219 -200 -1199 -199
rect -1546 -208 -1526 -207
rect -1546 -211 -1526 -210
rect -1219 -203 -1199 -202
rect -1219 -208 -1199 -207
rect -1219 -211 -1199 -210
rect -1546 -247 -1526 -246
rect -1546 -250 -1526 -249
rect -1440 -247 -1420 -246
rect -1546 -255 -1526 -254
rect -1674 -271 -1673 -261
rect -1671 -271 -1670 -261
rect -1623 -271 -1622 -261
rect -1620 -271 -1619 -261
rect -1546 -258 -1526 -257
rect -1440 -250 -1420 -249
rect -1440 -255 -1420 -254
rect -1440 -258 -1420 -257
rect -1219 -247 -1199 -246
rect -1219 -250 -1199 -249
rect -1113 -247 -1093 -246
rect -1219 -255 -1199 -254
rect -1346 -271 -1345 -261
rect -1343 -271 -1342 -261
rect -1296 -271 -1295 -261
rect -1293 -271 -1292 -261
rect -1219 -258 -1199 -257
rect -1113 -250 -1093 -249
rect -1113 -255 -1093 -254
rect -1113 -258 -1093 -257
rect -855 -294 -835 -293
rect -855 -297 -835 -296
rect -855 -302 -835 -301
rect -855 -305 -835 -304
rect -793 -325 -792 -315
rect -790 -325 -789 -315
rect -1440 -357 -1420 -356
rect -1440 -360 -1420 -359
rect -1113 -357 -1093 -356
rect -1440 -365 -1420 -364
rect -1440 -368 -1420 -367
rect -1113 -360 -1093 -359
rect -1113 -365 -1093 -364
rect -1546 -375 -1526 -374
rect -1546 -378 -1526 -377
rect -1113 -368 -1093 -367
rect -752 -370 -732 -369
rect -1219 -375 -1199 -374
rect -1546 -383 -1526 -382
rect -1546 -386 -1526 -385
rect -1219 -378 -1199 -377
rect -752 -373 -732 -372
rect -752 -378 -732 -377
rect -1219 -383 -1199 -382
rect -752 -381 -732 -380
rect -1219 -386 -1199 -385
rect -1546 -422 -1526 -421
rect -1546 -425 -1526 -424
rect -1440 -422 -1420 -421
rect -843 -404 -823 -403
rect -843 -407 -823 -406
rect -656 -404 -636 -403
rect -843 -412 -823 -411
rect -1546 -430 -1526 -429
rect -1674 -446 -1673 -436
rect -1671 -446 -1670 -436
rect -1623 -446 -1622 -436
rect -1620 -446 -1619 -436
rect -1546 -433 -1526 -432
rect -1440 -425 -1420 -424
rect -1440 -430 -1420 -429
rect -1440 -433 -1420 -432
rect -1219 -422 -1199 -421
rect -1219 -425 -1199 -424
rect -843 -415 -823 -414
rect -656 -407 -636 -406
rect -656 -412 -636 -411
rect -656 -415 -636 -414
rect -1113 -422 -1093 -421
rect -1219 -430 -1199 -429
rect -1346 -446 -1345 -436
rect -1343 -446 -1342 -436
rect -1296 -446 -1295 -436
rect -1293 -446 -1292 -436
rect -1219 -433 -1199 -432
rect -1113 -425 -1093 -424
rect -752 -426 -732 -425
rect -1113 -430 -1093 -429
rect -1113 -433 -1093 -432
rect -752 -429 -732 -428
rect -752 -434 -732 -433
rect -752 -437 -732 -436
<< pdiffusion >>
rect -1475 1529 -1455 1530
rect -1475 1526 -1455 1527
rect -1475 1521 -1455 1522
rect -1148 1529 -1128 1530
rect -1148 1526 -1128 1527
rect -1475 1518 -1455 1519
rect -1581 1511 -1561 1512
rect -1148 1521 -1128 1522
rect -1148 1518 -1128 1519
rect -1581 1508 -1561 1509
rect -1581 1503 -1561 1504
rect -1254 1511 -1234 1512
rect -1254 1508 -1234 1509
rect -1581 1500 -1561 1501
rect -1254 1503 -1234 1504
rect -1254 1500 -1234 1501
rect -400 1488 -399 1508
rect -397 1488 -396 1508
rect -1673 1464 -1672 1484
rect -1670 1464 -1669 1484
rect -1622 1464 -1621 1484
rect -1619 1464 -1618 1484
rect -1581 1464 -1561 1465
rect -1581 1461 -1561 1462
rect -1581 1456 -1561 1457
rect -1475 1464 -1455 1465
rect -1345 1464 -1344 1484
rect -1342 1464 -1341 1484
rect -1295 1464 -1294 1484
rect -1292 1464 -1291 1484
rect -477 1482 -457 1483
rect -477 1479 -457 1480
rect -477 1474 -457 1475
rect -477 1471 -457 1472
rect -1475 1461 -1455 1462
rect -1581 1453 -1561 1454
rect -1475 1456 -1455 1457
rect -1475 1453 -1455 1454
rect -1254 1464 -1234 1465
rect -1254 1461 -1234 1462
rect -1254 1456 -1234 1457
rect -1148 1464 -1128 1465
rect -1148 1461 -1128 1462
rect -1254 1453 -1234 1454
rect -1148 1456 -1128 1457
rect -1148 1453 -1128 1454
rect -252 1453 -251 1473
rect -249 1453 -248 1473
rect -339 1446 -299 1447
rect -339 1443 -299 1444
rect -339 1438 -299 1439
rect -339 1435 -299 1436
rect -887 1380 -867 1381
rect -887 1377 -867 1378
rect -887 1372 -867 1373
rect -789 1373 -788 1393
rect -786 1373 -785 1393
rect -887 1369 -867 1370
rect -57 1365 -37 1366
rect -57 1362 -37 1363
rect -1475 1351 -1455 1352
rect -1475 1348 -1455 1349
rect -1475 1343 -1455 1344
rect -1148 1351 -1128 1352
rect -57 1357 -37 1358
rect -57 1354 -37 1355
rect -1148 1348 -1128 1349
rect -1475 1340 -1455 1341
rect -1581 1333 -1561 1334
rect -1148 1343 -1128 1344
rect -1148 1340 -1128 1341
rect -1581 1330 -1561 1331
rect -1581 1325 -1561 1326
rect -1254 1333 -1234 1334
rect -1254 1330 -1234 1331
rect -1581 1322 -1561 1323
rect -1254 1325 -1234 1326
rect -148 1331 -128 1332
rect -148 1328 -128 1329
rect -1254 1322 -1234 1323
rect -148 1323 -128 1324
rect 39 1331 59 1332
rect 39 1328 59 1329
rect -148 1320 -128 1321
rect 39 1323 59 1324
rect 39 1320 59 1321
rect -1673 1286 -1672 1306
rect -1670 1286 -1669 1306
rect -1622 1286 -1621 1306
rect -1619 1286 -1618 1306
rect -1581 1286 -1561 1287
rect -1581 1283 -1561 1284
rect -1581 1278 -1561 1279
rect -1475 1286 -1455 1287
rect -1345 1286 -1344 1306
rect -1342 1286 -1341 1306
rect -1295 1286 -1294 1306
rect -1292 1286 -1291 1306
rect -784 1304 -764 1305
rect -57 1309 -37 1310
rect -57 1306 -37 1307
rect -784 1301 -764 1302
rect -784 1296 -764 1297
rect -57 1301 -37 1302
rect -57 1298 -37 1299
rect -784 1293 -764 1294
rect -1475 1283 -1455 1284
rect -1581 1275 -1561 1276
rect -1475 1278 -1455 1279
rect -1475 1275 -1455 1276
rect -1254 1286 -1234 1287
rect -1254 1283 -1234 1284
rect -1254 1278 -1234 1279
rect -1148 1286 -1128 1287
rect -1148 1283 -1128 1284
rect -1254 1275 -1234 1276
rect -1148 1278 -1128 1279
rect -1148 1275 -1128 1276
rect -875 1270 -855 1271
rect -875 1267 -855 1268
rect -875 1262 -855 1263
rect -688 1270 -668 1271
rect -688 1267 -668 1268
rect -875 1259 -855 1260
rect -688 1262 -668 1263
rect -688 1259 -668 1260
rect -784 1248 -764 1249
rect -784 1245 -764 1246
rect -784 1240 -764 1241
rect -784 1237 -764 1238
rect -488 1197 -468 1198
rect -488 1194 -468 1195
rect -488 1189 -468 1190
rect -402 1192 -401 1212
rect -399 1192 -398 1212
rect -29 1198 -9 1199
rect -29 1195 -9 1196
rect -488 1186 -468 1187
rect -1476 1176 -1456 1177
rect -1476 1173 -1456 1174
rect -1476 1168 -1456 1169
rect -1149 1176 -1129 1177
rect -488 1181 -468 1182
rect -488 1178 -468 1179
rect -29 1190 -9 1191
rect -29 1187 -9 1188
rect -1149 1173 -1129 1174
rect -1476 1165 -1456 1166
rect -1582 1158 -1562 1159
rect -1149 1168 -1129 1169
rect -1149 1165 -1129 1166
rect -1582 1155 -1562 1156
rect -1582 1150 -1562 1151
rect -1255 1158 -1235 1159
rect -120 1164 -100 1165
rect -120 1161 -100 1162
rect -1255 1155 -1235 1156
rect -1582 1147 -1562 1148
rect -1255 1150 -1235 1151
rect -120 1156 -100 1157
rect 67 1164 87 1165
rect 67 1161 87 1162
rect -120 1153 -100 1154
rect 67 1156 87 1157
rect 67 1153 87 1154
rect -1255 1147 -1235 1148
rect -29 1142 -9 1143
rect -29 1139 -9 1140
rect -1674 1111 -1673 1131
rect -1671 1111 -1670 1131
rect -1623 1111 -1622 1131
rect -1620 1111 -1619 1131
rect -1582 1111 -1562 1112
rect -1582 1108 -1562 1109
rect -1582 1103 -1562 1104
rect -1476 1111 -1456 1112
rect -1346 1111 -1345 1131
rect -1343 1111 -1342 1131
rect -1296 1111 -1295 1131
rect -1293 1111 -1292 1131
rect -404 1118 -403 1138
rect -401 1118 -400 1138
rect -29 1134 -9 1135
rect -29 1131 -9 1132
rect -1476 1108 -1456 1109
rect -1582 1100 -1562 1101
rect -1476 1103 -1456 1104
rect -1476 1100 -1456 1101
rect -1255 1111 -1235 1112
rect -1255 1108 -1235 1109
rect -1255 1103 -1235 1104
rect -1149 1111 -1129 1112
rect -481 1112 -461 1113
rect -481 1109 -461 1110
rect -1149 1108 -1129 1109
rect -1255 1100 -1235 1101
rect -1149 1103 -1129 1104
rect -481 1104 -461 1105
rect -481 1101 -461 1102
rect -1149 1100 -1129 1101
rect -292 1083 -232 1084
rect -292 1080 -232 1081
rect -292 1075 -232 1076
rect -186 1079 -185 1099
rect -183 1079 -182 1099
rect -292 1072 -232 1073
rect -292 1067 -232 1068
rect -292 1064 -232 1065
rect -891 1014 -871 1015
rect -891 1011 -871 1012
rect -1476 1001 -1456 1002
rect -1476 998 -1456 999
rect -1476 993 -1456 994
rect -1149 1001 -1129 1002
rect -891 1006 -871 1007
rect -793 1007 -792 1027
rect -790 1007 -789 1027
rect -891 1003 -871 1004
rect -1149 998 -1129 999
rect -1476 990 -1456 991
rect -1582 983 -1562 984
rect -1149 993 -1129 994
rect -1149 990 -1129 991
rect -1582 980 -1562 981
rect -1582 975 -1562 976
rect -1255 983 -1235 984
rect -1255 980 -1235 981
rect -1582 972 -1562 973
rect -1255 975 -1235 976
rect -1255 972 -1235 973
rect -1674 936 -1673 956
rect -1671 936 -1670 956
rect -1623 936 -1622 956
rect -1620 936 -1619 956
rect -1582 936 -1562 937
rect -1582 933 -1562 934
rect -1582 928 -1562 929
rect -1476 936 -1456 937
rect -1346 936 -1345 956
rect -1343 936 -1342 956
rect -1296 936 -1295 956
rect -1293 936 -1292 956
rect -1476 933 -1456 934
rect -1582 925 -1562 926
rect -1476 928 -1456 929
rect -1476 925 -1456 926
rect -1255 936 -1235 937
rect -1255 933 -1235 934
rect -1255 928 -1235 929
rect -1149 936 -1129 937
rect -788 938 -768 939
rect -788 935 -768 936
rect -1149 933 -1129 934
rect -1255 925 -1235 926
rect -1149 928 -1129 929
rect -788 930 -768 931
rect -788 927 -768 928
rect -1149 925 -1129 926
rect -879 904 -859 905
rect -879 901 -859 902
rect -879 896 -859 897
rect -692 904 -672 905
rect -692 901 -672 902
rect -879 893 -859 894
rect -692 896 -672 897
rect -692 893 -672 894
rect -788 882 -768 883
rect -788 879 -768 880
rect -788 874 -768 875
rect 79 879 99 880
rect 79 876 99 877
rect -788 871 -768 872
rect 79 871 99 872
rect 79 868 99 869
rect -448 847 -428 848
rect -448 844 -428 845
rect -448 839 -428 840
rect -352 839 -351 859
rect -349 839 -348 859
rect -227 846 -147 847
rect -227 843 -147 844
rect -448 836 -428 837
rect -1476 825 -1456 826
rect -1476 822 -1456 823
rect -1476 817 -1456 818
rect -1149 825 -1129 826
rect -448 831 -428 832
rect -448 828 -428 829
rect -1149 822 -1129 823
rect -1476 814 -1456 815
rect -1582 807 -1562 808
rect -1149 817 -1129 818
rect -448 823 -428 824
rect -227 838 -147 839
rect -100 836 -99 856
rect -97 836 -96 856
rect -12 845 8 846
rect -12 842 8 843
rect -227 835 -147 836
rect -227 830 -147 831
rect -227 827 -147 828
rect -448 820 -428 821
rect -1149 814 -1129 815
rect -1582 804 -1562 805
rect -1582 799 -1562 800
rect -1255 807 -1235 808
rect -227 822 -147 823
rect -12 837 8 838
rect 175 845 195 846
rect 175 842 195 843
rect -12 834 8 835
rect 175 837 195 838
rect 175 834 195 835
rect 79 823 99 824
rect 79 820 99 821
rect -227 819 -147 820
rect 79 815 99 816
rect 79 812 99 813
rect -1255 804 -1235 805
rect -1582 796 -1562 797
rect -1255 799 -1235 800
rect -1255 796 -1235 797
rect -1674 760 -1673 780
rect -1671 760 -1670 780
rect -1623 760 -1622 780
rect -1620 760 -1619 780
rect -1582 760 -1562 761
rect -1582 757 -1562 758
rect -1582 752 -1562 753
rect -1476 760 -1456 761
rect -1346 760 -1345 780
rect -1343 760 -1342 780
rect -1296 760 -1295 780
rect -1293 760 -1292 780
rect -446 774 -426 775
rect -446 771 -426 772
rect -1476 757 -1456 758
rect -1582 749 -1562 750
rect -1476 752 -1456 753
rect -1476 749 -1456 750
rect -1255 760 -1235 761
rect -1255 757 -1235 758
rect -1255 752 -1235 753
rect -1149 760 -1129 761
rect -446 766 -426 767
rect -360 769 -359 789
rect -357 769 -356 789
rect -446 763 -426 764
rect -1149 757 -1129 758
rect -1255 749 -1235 750
rect -1149 752 -1129 753
rect -446 758 -426 759
rect -446 755 -426 756
rect -1149 749 -1129 750
rect -369 694 -368 714
rect -366 694 -365 714
rect -446 688 -426 689
rect -446 685 -426 686
rect -446 680 -426 681
rect -446 677 -426 678
rect -1476 650 -1456 651
rect -1476 647 -1456 648
rect -1476 642 -1456 643
rect -1149 650 -1129 651
rect -891 656 -871 657
rect -891 653 -871 654
rect -1149 647 -1129 648
rect -1476 639 -1456 640
rect -1582 632 -1562 633
rect -1149 642 -1129 643
rect -891 648 -871 649
rect -793 649 -792 669
rect -790 649 -789 669
rect -891 645 -871 646
rect -1149 639 -1129 640
rect -1582 629 -1562 630
rect -1582 624 -1562 625
rect -1255 632 -1235 633
rect -1255 629 -1235 630
rect -1582 621 -1562 622
rect -1255 624 -1235 625
rect -1255 621 -1235 622
rect -1674 585 -1673 605
rect -1671 585 -1670 605
rect -1623 585 -1622 605
rect -1620 585 -1619 605
rect -1582 585 -1562 586
rect -1582 582 -1562 583
rect -1582 577 -1562 578
rect -1476 585 -1456 586
rect -1346 585 -1345 605
rect -1343 585 -1342 605
rect -1296 585 -1295 605
rect -1293 585 -1292 605
rect -1476 582 -1456 583
rect -1582 574 -1562 575
rect -1476 577 -1456 578
rect -1476 574 -1456 575
rect -1255 585 -1235 586
rect -1255 582 -1235 583
rect -1255 577 -1235 578
rect -1149 585 -1129 586
rect -1149 582 -1129 583
rect -1255 574 -1235 575
rect -1149 577 -1129 578
rect -788 580 -768 581
rect -788 577 -768 578
rect -1149 574 -1129 575
rect -788 572 -768 573
rect -788 569 -768 570
rect -879 546 -859 547
rect -879 543 -859 544
rect -879 538 -859 539
rect -692 546 -672 547
rect -692 543 -672 544
rect -879 535 -859 536
rect -692 538 -672 539
rect -692 535 -672 536
rect -788 524 -768 525
rect -788 521 -768 522
rect -788 516 -768 517
rect -788 513 -768 514
rect -1475 344 -1455 345
rect -1475 341 -1455 342
rect -1475 336 -1455 337
rect -1148 344 -1128 345
rect -1148 341 -1128 342
rect -1475 333 -1455 334
rect -1581 326 -1561 327
rect -1148 336 -1128 337
rect -1148 333 -1128 334
rect -1581 323 -1561 324
rect -1581 318 -1561 319
rect -1254 326 -1234 327
rect -1254 323 -1234 324
rect -1581 315 -1561 316
rect -1254 318 -1234 319
rect -1254 315 -1234 316
rect -1673 279 -1672 299
rect -1670 279 -1669 299
rect -1622 279 -1621 299
rect -1619 279 -1618 299
rect -1581 279 -1561 280
rect -1581 276 -1561 277
rect -1581 271 -1561 272
rect -1475 279 -1455 280
rect -1345 279 -1344 299
rect -1342 279 -1341 299
rect -1295 279 -1294 299
rect -1292 279 -1291 299
rect -1475 276 -1455 277
rect -1581 268 -1561 269
rect -1475 271 -1455 272
rect -1475 268 -1455 269
rect -1254 279 -1234 280
rect -1254 276 -1234 277
rect -1254 271 -1234 272
rect -1148 279 -1128 280
rect -1148 276 -1128 277
rect -1254 268 -1234 269
rect -1148 271 -1128 272
rect -1148 268 -1128 269
rect -891 209 -871 210
rect -891 206 -871 207
rect -891 201 -871 202
rect -793 202 -792 222
rect -790 202 -789 222
rect -891 198 -871 199
rect -1476 169 -1456 170
rect -1476 166 -1456 167
rect -1476 161 -1456 162
rect -1149 169 -1129 170
rect -1149 166 -1129 167
rect -1476 158 -1456 159
rect -1582 151 -1562 152
rect -1149 161 -1129 162
rect -1149 158 -1129 159
rect -1582 148 -1562 149
rect -1582 143 -1562 144
rect -1255 151 -1235 152
rect -1255 148 -1235 149
rect -1582 140 -1562 141
rect -1255 143 -1235 144
rect -1255 140 -1235 141
rect -788 133 -768 134
rect -788 130 -768 131
rect -1674 104 -1673 124
rect -1671 104 -1670 124
rect -1623 104 -1622 124
rect -1620 104 -1619 124
rect -1582 104 -1562 105
rect -1582 101 -1562 102
rect -1582 96 -1562 97
rect -1476 104 -1456 105
rect -1346 104 -1345 124
rect -1343 104 -1342 124
rect -1296 104 -1295 124
rect -1293 104 -1292 124
rect -788 125 -768 126
rect -788 122 -768 123
rect -1476 101 -1456 102
rect -1582 93 -1562 94
rect -1476 96 -1456 97
rect -1476 93 -1456 94
rect -1255 104 -1235 105
rect -1255 101 -1235 102
rect -1255 96 -1235 97
rect -1149 104 -1129 105
rect -1149 101 -1129 102
rect -1255 93 -1235 94
rect -1149 96 -1129 97
rect -879 99 -859 100
rect -879 96 -859 97
rect -1149 93 -1129 94
rect -879 91 -859 92
rect -692 99 -672 100
rect -692 96 -672 97
rect -879 88 -859 89
rect -692 91 -672 92
rect -692 88 -672 89
rect -788 77 -768 78
rect -788 74 -768 75
rect -788 69 -768 70
rect -788 66 -768 67
rect -1476 -6 -1456 -5
rect -1476 -9 -1456 -8
rect -1476 -14 -1456 -13
rect -1149 -6 -1129 -5
rect -1149 -9 -1129 -8
rect -1476 -17 -1456 -16
rect -1582 -24 -1562 -23
rect -1149 -14 -1129 -13
rect -1149 -17 -1129 -16
rect -1582 -27 -1562 -26
rect -1582 -32 -1562 -31
rect -1255 -24 -1235 -23
rect -1255 -27 -1235 -26
rect -1582 -35 -1562 -34
rect -1255 -32 -1235 -31
rect -1255 -35 -1235 -34
rect -1674 -71 -1673 -51
rect -1671 -71 -1670 -51
rect -1623 -71 -1622 -51
rect -1620 -71 -1619 -51
rect -1582 -71 -1562 -70
rect -1582 -74 -1562 -73
rect -1582 -79 -1562 -78
rect -1476 -71 -1456 -70
rect -1346 -71 -1345 -51
rect -1343 -71 -1342 -51
rect -1296 -71 -1295 -51
rect -1293 -71 -1292 -51
rect -1476 -74 -1456 -73
rect -1582 -82 -1562 -81
rect -1476 -79 -1456 -78
rect -1476 -82 -1456 -81
rect -1255 -71 -1235 -70
rect -1255 -74 -1235 -73
rect -1255 -79 -1235 -78
rect -1149 -71 -1129 -70
rect -1149 -74 -1129 -73
rect -1255 -82 -1235 -81
rect -1149 -79 -1129 -78
rect -1149 -82 -1129 -81
rect -1476 -182 -1456 -181
rect -1476 -185 -1456 -184
rect -1476 -190 -1456 -189
rect -1149 -182 -1129 -181
rect -1149 -185 -1129 -184
rect -1476 -193 -1456 -192
rect -1582 -200 -1562 -199
rect -1149 -190 -1129 -189
rect -1149 -193 -1129 -192
rect -1582 -203 -1562 -202
rect -1582 -208 -1562 -207
rect -1255 -200 -1235 -199
rect -1255 -203 -1235 -202
rect -1582 -211 -1562 -210
rect -1255 -208 -1235 -207
rect -1255 -211 -1235 -210
rect -1674 -247 -1673 -227
rect -1671 -247 -1670 -227
rect -1623 -247 -1622 -227
rect -1620 -247 -1619 -227
rect -1582 -247 -1562 -246
rect -1582 -250 -1562 -249
rect -1582 -255 -1562 -254
rect -1476 -247 -1456 -246
rect -1346 -247 -1345 -227
rect -1343 -247 -1342 -227
rect -1296 -247 -1295 -227
rect -1293 -247 -1292 -227
rect -1476 -250 -1456 -249
rect -1582 -258 -1562 -257
rect -1476 -255 -1456 -254
rect -1476 -258 -1456 -257
rect -1255 -247 -1235 -246
rect -1255 -250 -1235 -249
rect -1255 -255 -1235 -254
rect -1149 -247 -1129 -246
rect -1149 -250 -1129 -249
rect -1255 -258 -1235 -257
rect -1149 -255 -1129 -254
rect -1149 -258 -1129 -257
rect -891 -294 -871 -293
rect -891 -297 -871 -296
rect -891 -302 -871 -301
rect -793 -301 -792 -281
rect -790 -301 -789 -281
rect -891 -305 -871 -304
rect -1476 -357 -1456 -356
rect -1476 -360 -1456 -359
rect -1476 -365 -1456 -364
rect -1149 -357 -1129 -356
rect -1149 -360 -1129 -359
rect -1476 -368 -1456 -367
rect -1582 -375 -1562 -374
rect -1149 -365 -1129 -364
rect -1149 -368 -1129 -367
rect -1582 -378 -1562 -377
rect -1582 -383 -1562 -382
rect -1255 -375 -1235 -374
rect -788 -370 -768 -369
rect -788 -373 -768 -372
rect -1255 -378 -1235 -377
rect -1582 -386 -1562 -385
rect -1255 -383 -1235 -382
rect -788 -378 -768 -377
rect -788 -381 -768 -380
rect -1255 -386 -1235 -385
rect -1674 -422 -1673 -402
rect -1671 -422 -1670 -402
rect -1623 -422 -1622 -402
rect -1620 -422 -1619 -402
rect -1582 -422 -1562 -421
rect -1582 -425 -1562 -424
rect -1582 -430 -1562 -429
rect -1476 -422 -1456 -421
rect -1346 -422 -1345 -402
rect -1343 -422 -1342 -402
rect -1296 -422 -1295 -402
rect -1293 -422 -1292 -402
rect -879 -404 -859 -403
rect -879 -407 -859 -406
rect -879 -412 -859 -411
rect -692 -404 -672 -403
rect -692 -407 -672 -406
rect -879 -415 -859 -414
rect -1476 -425 -1456 -424
rect -1582 -433 -1562 -432
rect -1476 -430 -1456 -429
rect -1476 -433 -1456 -432
rect -1255 -422 -1235 -421
rect -1255 -425 -1235 -424
rect -1255 -430 -1235 -429
rect -1149 -422 -1129 -421
rect -692 -412 -672 -411
rect -692 -415 -672 -414
rect -1149 -425 -1129 -424
rect -1255 -433 -1235 -432
rect -1149 -430 -1129 -429
rect -788 -426 -768 -425
rect -788 -429 -768 -428
rect -1149 -433 -1129 -432
rect -788 -434 -768 -433
rect -788 -437 -768 -436
<< ndcontact >>
rect -1439 1530 -1419 1534
rect -1112 1530 -1092 1534
rect -1439 1522 -1419 1526
rect -1545 1512 -1525 1516
rect -1112 1522 -1092 1526
rect -1439 1514 -1419 1518
rect -1218 1512 -1198 1516
rect -1112 1514 -1092 1518
rect -1545 1504 -1525 1508
rect -1218 1504 -1198 1508
rect -1545 1496 -1525 1500
rect -1218 1496 -1198 1500
rect -1545 1465 -1525 1469
rect -1439 1465 -1419 1469
rect -444 1483 -424 1487
rect -444 1475 -424 1479
rect -1545 1457 -1525 1461
rect -1677 1440 -1673 1450
rect -1669 1440 -1665 1450
rect -1626 1440 -1622 1450
rect -1618 1440 -1614 1450
rect -1439 1457 -1419 1461
rect -1545 1449 -1525 1453
rect -1439 1449 -1419 1453
rect -1218 1465 -1198 1469
rect -1112 1465 -1092 1469
rect -444 1467 -424 1471
rect -404 1462 -400 1472
rect -396 1462 -392 1472
rect -1218 1457 -1198 1461
rect -1349 1440 -1345 1450
rect -1341 1440 -1337 1450
rect -1299 1440 -1295 1450
rect -1291 1440 -1287 1450
rect -1112 1457 -1092 1461
rect -1218 1449 -1198 1453
rect -1112 1449 -1092 1453
rect -287 1447 -277 1451
rect -287 1439 -277 1443
rect -287 1431 -277 1435
rect -256 1427 -252 1437
rect -248 1427 -244 1437
rect -851 1381 -831 1385
rect -851 1373 -831 1377
rect -851 1365 -831 1369
rect -21 1366 -1 1370
rect -1439 1352 -1419 1356
rect -1112 1352 -1092 1356
rect -793 1349 -789 1359
rect -785 1349 -781 1359
rect -21 1358 -1 1362
rect -21 1350 -1 1354
rect -1439 1344 -1419 1348
rect -1545 1334 -1525 1338
rect -1112 1344 -1092 1348
rect -1439 1336 -1419 1340
rect -1218 1334 -1198 1338
rect -1112 1336 -1092 1340
rect -1545 1326 -1525 1330
rect -1218 1326 -1198 1330
rect -112 1332 -92 1336
rect -1545 1318 -1525 1322
rect -1218 1318 -1198 1322
rect 75 1332 95 1336
rect -112 1324 -92 1328
rect 75 1324 95 1328
rect -112 1316 -92 1320
rect 75 1316 95 1320
rect -1545 1287 -1525 1291
rect -1439 1287 -1419 1291
rect -748 1305 -728 1309
rect -21 1310 -1 1314
rect -748 1297 -728 1301
rect -21 1302 -1 1306
rect -21 1294 -1 1298
rect -1545 1279 -1525 1283
rect -1677 1262 -1673 1272
rect -1669 1262 -1665 1272
rect -1626 1262 -1622 1272
rect -1618 1262 -1614 1272
rect -1439 1279 -1419 1283
rect -1545 1271 -1525 1275
rect -1439 1271 -1419 1275
rect -1218 1287 -1198 1291
rect -1112 1287 -1092 1291
rect -748 1289 -728 1293
rect -1218 1279 -1198 1283
rect -1349 1262 -1345 1272
rect -1341 1262 -1337 1272
rect -1299 1262 -1295 1272
rect -1291 1262 -1287 1272
rect -1112 1279 -1092 1283
rect -1218 1271 -1198 1275
rect -1112 1271 -1092 1275
rect -839 1271 -819 1275
rect -652 1271 -632 1275
rect -839 1263 -819 1267
rect -652 1263 -632 1267
rect -839 1255 -819 1259
rect -652 1255 -632 1259
rect -748 1249 -728 1253
rect -748 1241 -728 1245
rect -748 1233 -728 1237
rect -456 1198 -426 1202
rect -456 1190 -426 1194
rect 7 1199 27 1203
rect -1440 1177 -1420 1181
rect -1113 1177 -1093 1181
rect -456 1182 -426 1186
rect -456 1174 -426 1178
rect 7 1191 27 1195
rect 7 1183 27 1187
rect -1440 1169 -1420 1173
rect -1546 1159 -1526 1163
rect -1113 1169 -1093 1173
rect -406 1166 -402 1176
rect -398 1166 -394 1176
rect -1440 1161 -1420 1165
rect -1219 1159 -1199 1163
rect -1113 1161 -1093 1165
rect -84 1165 -64 1169
rect -1546 1151 -1526 1155
rect -1219 1151 -1199 1155
rect 103 1165 123 1169
rect -84 1157 -64 1161
rect 103 1157 123 1161
rect -84 1149 -64 1153
rect 103 1149 123 1153
rect -1546 1143 -1526 1147
rect -1219 1143 -1199 1147
rect 7 1143 27 1147
rect -1546 1112 -1526 1116
rect -1440 1112 -1420 1116
rect 7 1135 27 1139
rect 7 1127 27 1131
rect -1546 1104 -1526 1108
rect -1678 1087 -1674 1097
rect -1670 1087 -1666 1097
rect -1627 1087 -1623 1097
rect -1619 1087 -1615 1097
rect -1440 1104 -1420 1108
rect -1546 1096 -1526 1100
rect -1440 1096 -1420 1100
rect -1219 1112 -1199 1116
rect -1113 1112 -1093 1116
rect -448 1113 -428 1117
rect -1219 1104 -1199 1108
rect -1350 1087 -1346 1097
rect -1342 1087 -1338 1097
rect -1300 1087 -1296 1097
rect -1292 1087 -1288 1097
rect -1113 1104 -1093 1108
rect -448 1105 -428 1109
rect -1219 1096 -1199 1100
rect -1113 1096 -1093 1100
rect -448 1097 -428 1101
rect -408 1092 -404 1102
rect -400 1092 -396 1102
rect -220 1084 -210 1088
rect -220 1076 -210 1080
rect -220 1068 -210 1072
rect -220 1060 -210 1064
rect -190 1053 -186 1063
rect -182 1053 -178 1063
rect -855 1015 -835 1019
rect -1440 1002 -1420 1006
rect -1113 1002 -1093 1006
rect -855 1007 -835 1011
rect -855 999 -835 1003
rect -1440 994 -1420 998
rect -1546 984 -1526 988
rect -1113 994 -1093 998
rect -1440 986 -1420 990
rect -1219 984 -1199 988
rect -1113 986 -1093 990
rect -797 983 -793 993
rect -789 983 -785 993
rect -1546 976 -1526 980
rect -1219 976 -1199 980
rect -1546 968 -1526 972
rect -1219 968 -1199 972
rect -1546 937 -1526 941
rect -1440 937 -1420 941
rect -1546 929 -1526 933
rect -1678 912 -1674 922
rect -1670 912 -1666 922
rect -1627 912 -1623 922
rect -1619 912 -1615 922
rect -1440 929 -1420 933
rect -1546 921 -1526 925
rect -1440 921 -1420 925
rect -1219 937 -1199 941
rect -1113 937 -1093 941
rect -752 939 -732 943
rect -1219 929 -1199 933
rect -1350 912 -1346 922
rect -1342 912 -1338 922
rect -1300 912 -1296 922
rect -1292 912 -1288 922
rect -1113 929 -1093 933
rect -752 931 -732 935
rect -1219 921 -1199 925
rect -1113 921 -1093 925
rect -752 923 -732 927
rect -843 905 -823 909
rect -656 905 -636 909
rect -843 897 -823 901
rect -656 897 -636 901
rect -843 889 -823 893
rect -656 889 -636 893
rect -752 883 -732 887
rect -752 875 -732 879
rect 115 880 135 884
rect -752 867 -732 871
rect 115 872 135 876
rect 115 864 135 868
rect -416 848 -376 852
rect -416 840 -376 844
rect -135 847 -125 851
rect -1440 826 -1420 830
rect -1113 826 -1093 830
rect -416 832 -376 836
rect -1440 818 -1420 822
rect -1546 808 -1526 812
rect -1113 818 -1093 822
rect -416 824 -376 828
rect -135 839 -125 843
rect 24 846 44 850
rect -135 831 -125 835
rect -416 816 -376 820
rect -1440 810 -1420 814
rect -1219 808 -1199 812
rect -1113 810 -1093 814
rect -356 813 -352 823
rect -348 813 -344 823
rect -135 823 -125 827
rect 211 846 231 850
rect 24 838 44 842
rect 211 838 231 842
rect 24 830 44 834
rect 211 830 231 834
rect 115 824 135 828
rect -135 815 -125 819
rect -104 810 -100 820
rect -96 810 -92 820
rect 115 816 135 820
rect 115 808 135 812
rect -1546 800 -1526 804
rect -1219 800 -1199 804
rect -1546 792 -1526 796
rect -1219 792 -1199 796
rect -1546 761 -1526 765
rect -1440 761 -1420 765
rect -414 775 -384 779
rect -1546 753 -1526 757
rect -1678 736 -1674 746
rect -1670 736 -1666 746
rect -1627 736 -1623 746
rect -1619 736 -1615 746
rect -1440 753 -1420 757
rect -1546 745 -1526 749
rect -1440 745 -1420 749
rect -1219 761 -1199 765
rect -1113 761 -1093 765
rect -414 767 -384 771
rect -1219 753 -1199 757
rect -1350 736 -1346 746
rect -1342 736 -1338 746
rect -1300 736 -1296 746
rect -1292 736 -1288 746
rect -1113 753 -1093 757
rect -414 759 -384 763
rect -414 751 -384 755
rect -1219 745 -1199 749
rect -1113 745 -1093 749
rect -364 743 -360 753
rect -356 743 -352 753
rect -413 689 -393 693
rect -413 681 -393 685
rect -413 673 -393 677
rect -1440 651 -1420 655
rect -1113 651 -1093 655
rect -855 657 -835 661
rect -1440 643 -1420 647
rect -1546 633 -1526 637
rect -1113 643 -1093 647
rect -855 649 -835 653
rect -373 668 -369 678
rect -365 668 -361 678
rect -855 641 -835 645
rect -1440 635 -1420 639
rect -1219 633 -1199 637
rect -1113 635 -1093 639
rect -1546 625 -1526 629
rect -1219 625 -1199 629
rect -797 625 -793 635
rect -789 625 -785 635
rect -1546 617 -1526 621
rect -1219 617 -1199 621
rect -1546 586 -1526 590
rect -1440 586 -1420 590
rect -1546 578 -1526 582
rect -1678 561 -1674 571
rect -1670 561 -1666 571
rect -1627 561 -1623 571
rect -1619 561 -1615 571
rect -1440 578 -1420 582
rect -1546 570 -1526 574
rect -1440 570 -1420 574
rect -1219 586 -1199 590
rect -1113 586 -1093 590
rect -1219 578 -1199 582
rect -1350 561 -1346 571
rect -1342 561 -1338 571
rect -1300 561 -1296 571
rect -1292 561 -1288 571
rect -1113 578 -1093 582
rect -752 581 -732 585
rect -1219 570 -1199 574
rect -1113 570 -1093 574
rect -752 573 -732 577
rect -752 565 -732 569
rect -843 547 -823 551
rect -656 547 -636 551
rect -843 539 -823 543
rect -656 539 -636 543
rect -843 531 -823 535
rect -656 531 -636 535
rect -752 525 -732 529
rect -752 517 -732 521
rect -752 509 -732 513
rect -1439 345 -1419 349
rect -1112 345 -1092 349
rect -1439 337 -1419 341
rect -1545 327 -1525 331
rect -1112 337 -1092 341
rect -1439 329 -1419 333
rect -1218 327 -1198 331
rect -1112 329 -1092 333
rect -1545 319 -1525 323
rect -1218 319 -1198 323
rect -1545 311 -1525 315
rect -1218 311 -1198 315
rect -1545 280 -1525 284
rect -1439 280 -1419 284
rect -1545 272 -1525 276
rect -1677 255 -1673 265
rect -1669 255 -1665 265
rect -1626 255 -1622 265
rect -1618 255 -1614 265
rect -1439 272 -1419 276
rect -1545 264 -1525 268
rect -1439 264 -1419 268
rect -1218 280 -1198 284
rect -1112 280 -1092 284
rect -1218 272 -1198 276
rect -1349 255 -1345 265
rect -1341 255 -1337 265
rect -1299 255 -1295 265
rect -1291 255 -1287 265
rect -1112 272 -1092 276
rect -1218 264 -1198 268
rect -1112 264 -1092 268
rect -855 210 -835 214
rect -855 202 -835 206
rect -855 194 -835 198
rect -797 178 -793 188
rect -789 178 -785 188
rect -1440 170 -1420 174
rect -1113 170 -1093 174
rect -1440 162 -1420 166
rect -1546 152 -1526 156
rect -1113 162 -1093 166
rect -1440 154 -1420 158
rect -1219 152 -1199 156
rect -1113 154 -1093 158
rect -1546 144 -1526 148
rect -1219 144 -1199 148
rect -1546 136 -1526 140
rect -1219 136 -1199 140
rect -752 134 -732 138
rect -1546 105 -1526 109
rect -1440 105 -1420 109
rect -752 126 -732 130
rect -752 118 -732 122
rect -1546 97 -1526 101
rect -1678 80 -1674 90
rect -1670 80 -1666 90
rect -1627 80 -1623 90
rect -1619 80 -1615 90
rect -1440 97 -1420 101
rect -1546 89 -1526 93
rect -1440 89 -1420 93
rect -1219 105 -1199 109
rect -1113 105 -1093 109
rect -1219 97 -1199 101
rect -1350 80 -1346 90
rect -1342 80 -1338 90
rect -1300 80 -1296 90
rect -1292 80 -1288 90
rect -1113 97 -1093 101
rect -843 100 -823 104
rect -1219 89 -1199 93
rect -1113 89 -1093 93
rect -656 100 -636 104
rect -843 92 -823 96
rect -656 92 -636 96
rect -843 84 -823 88
rect -656 84 -636 88
rect -752 78 -732 82
rect -752 70 -732 74
rect -752 62 -732 66
rect -1440 -5 -1420 -1
rect -1113 -5 -1093 -1
rect -1440 -13 -1420 -9
rect -1546 -23 -1526 -19
rect -1113 -13 -1093 -9
rect -1440 -21 -1420 -17
rect -1219 -23 -1199 -19
rect -1113 -21 -1093 -17
rect -1546 -31 -1526 -27
rect -1219 -31 -1199 -27
rect -1546 -39 -1526 -35
rect -1219 -39 -1199 -35
rect -1546 -70 -1526 -66
rect -1440 -70 -1420 -66
rect -1546 -78 -1526 -74
rect -1678 -95 -1674 -85
rect -1670 -95 -1666 -85
rect -1627 -95 -1623 -85
rect -1619 -95 -1615 -85
rect -1440 -78 -1420 -74
rect -1546 -86 -1526 -82
rect -1440 -86 -1420 -82
rect -1219 -70 -1199 -66
rect -1113 -70 -1093 -66
rect -1219 -78 -1199 -74
rect -1350 -95 -1346 -85
rect -1342 -95 -1338 -85
rect -1300 -95 -1296 -85
rect -1292 -95 -1288 -85
rect -1113 -78 -1093 -74
rect -1219 -86 -1199 -82
rect -1113 -86 -1093 -82
rect -1440 -181 -1420 -177
rect -1113 -181 -1093 -177
rect -1440 -189 -1420 -185
rect -1546 -199 -1526 -195
rect -1113 -189 -1093 -185
rect -1440 -197 -1420 -193
rect -1219 -199 -1199 -195
rect -1113 -197 -1093 -193
rect -1546 -207 -1526 -203
rect -1219 -207 -1199 -203
rect -1546 -215 -1526 -211
rect -1219 -215 -1199 -211
rect -1546 -246 -1526 -242
rect -1440 -246 -1420 -242
rect -1546 -254 -1526 -250
rect -1678 -271 -1674 -261
rect -1670 -271 -1666 -261
rect -1627 -271 -1623 -261
rect -1619 -271 -1615 -261
rect -1440 -254 -1420 -250
rect -1546 -262 -1526 -258
rect -1440 -262 -1420 -258
rect -1219 -246 -1199 -242
rect -1113 -246 -1093 -242
rect -1219 -254 -1199 -250
rect -1350 -271 -1346 -261
rect -1342 -271 -1338 -261
rect -1300 -271 -1296 -261
rect -1292 -271 -1288 -261
rect -1113 -254 -1093 -250
rect -1219 -262 -1199 -258
rect -1113 -262 -1093 -258
rect -855 -293 -835 -289
rect -855 -301 -835 -297
rect -855 -309 -835 -305
rect -797 -325 -793 -315
rect -789 -325 -785 -315
rect -1440 -356 -1420 -352
rect -1113 -356 -1093 -352
rect -1440 -364 -1420 -360
rect -1546 -374 -1526 -370
rect -1113 -364 -1093 -360
rect -1440 -372 -1420 -368
rect -1219 -374 -1199 -370
rect -1113 -372 -1093 -368
rect -752 -369 -732 -365
rect -1546 -382 -1526 -378
rect -1219 -382 -1199 -378
rect -752 -377 -732 -373
rect -752 -385 -732 -381
rect -1546 -390 -1526 -386
rect -1219 -390 -1199 -386
rect -1546 -421 -1526 -417
rect -1440 -421 -1420 -417
rect -843 -403 -823 -399
rect -656 -403 -636 -399
rect -843 -411 -823 -407
rect -1546 -429 -1526 -425
rect -1678 -446 -1674 -436
rect -1670 -446 -1666 -436
rect -1627 -446 -1623 -436
rect -1619 -446 -1615 -436
rect -1440 -429 -1420 -425
rect -1546 -437 -1526 -433
rect -1440 -437 -1420 -433
rect -1219 -421 -1199 -417
rect -1113 -421 -1093 -417
rect -656 -411 -636 -407
rect -843 -419 -823 -415
rect -656 -419 -636 -415
rect -1219 -429 -1199 -425
rect -1350 -446 -1346 -436
rect -1342 -446 -1338 -436
rect -1300 -446 -1296 -436
rect -1292 -446 -1288 -436
rect -1113 -429 -1093 -425
rect -752 -425 -732 -421
rect -1219 -437 -1199 -433
rect -1113 -437 -1093 -433
rect -752 -433 -732 -429
rect -752 -441 -732 -437
<< pdcontact >>
rect -1475 1530 -1455 1534
rect -1148 1530 -1128 1534
rect -1475 1522 -1455 1526
rect -1148 1522 -1128 1526
rect -1581 1512 -1561 1516
rect -1475 1514 -1455 1518
rect -1254 1512 -1234 1516
rect -1581 1504 -1561 1508
rect -1148 1514 -1128 1518
rect -1254 1504 -1234 1508
rect -1581 1496 -1561 1500
rect -1254 1496 -1234 1500
rect -404 1488 -400 1508
rect -396 1488 -392 1508
rect -1677 1464 -1673 1484
rect -1669 1464 -1665 1484
rect -1626 1464 -1622 1484
rect -1618 1464 -1614 1484
rect -1581 1465 -1561 1469
rect -1475 1465 -1455 1469
rect -1581 1457 -1561 1461
rect -1349 1464 -1345 1484
rect -1341 1464 -1337 1484
rect -1299 1464 -1295 1484
rect -1291 1464 -1287 1484
rect -477 1483 -457 1487
rect -477 1475 -457 1479
rect -1254 1465 -1234 1469
rect -1475 1457 -1455 1461
rect -1581 1449 -1561 1453
rect -1475 1449 -1455 1453
rect -1148 1465 -1128 1469
rect -1254 1457 -1234 1461
rect -477 1467 -457 1471
rect -1148 1457 -1128 1461
rect -1254 1449 -1234 1453
rect -1148 1449 -1128 1453
rect -256 1453 -252 1473
rect -248 1453 -244 1473
rect -339 1447 -299 1451
rect -339 1439 -299 1443
rect -339 1431 -299 1435
rect -887 1381 -867 1385
rect -887 1373 -867 1377
rect -793 1373 -789 1393
rect -785 1373 -781 1393
rect -887 1365 -867 1369
rect -57 1366 -37 1370
rect -1475 1352 -1455 1356
rect -1148 1352 -1128 1356
rect -1475 1344 -1455 1348
rect -57 1358 -37 1362
rect -57 1350 -37 1354
rect -1148 1344 -1128 1348
rect -1581 1334 -1561 1338
rect -1475 1336 -1455 1340
rect -1254 1334 -1234 1338
rect -1581 1326 -1561 1330
rect -1148 1336 -1128 1340
rect -148 1332 -128 1336
rect -1254 1326 -1234 1330
rect -1581 1318 -1561 1322
rect 39 1332 59 1336
rect -148 1324 -128 1328
rect -1254 1318 -1234 1322
rect 39 1324 59 1328
rect -148 1316 -128 1320
rect 39 1316 59 1320
rect -57 1310 -37 1314
rect -1677 1286 -1673 1306
rect -1669 1286 -1665 1306
rect -1626 1286 -1622 1306
rect -1618 1286 -1614 1306
rect -1581 1287 -1561 1291
rect -1475 1287 -1455 1291
rect -1581 1279 -1561 1283
rect -1349 1286 -1345 1306
rect -1341 1286 -1337 1306
rect -1299 1286 -1295 1306
rect -1291 1286 -1287 1306
rect -784 1305 -764 1309
rect -57 1302 -37 1306
rect -784 1297 -764 1301
rect -57 1294 -37 1298
rect -1254 1287 -1234 1291
rect -1475 1279 -1455 1283
rect -1581 1271 -1561 1275
rect -1475 1271 -1455 1275
rect -1148 1287 -1128 1291
rect -1254 1279 -1234 1283
rect -784 1289 -764 1293
rect -1148 1279 -1128 1283
rect -1254 1271 -1234 1275
rect -1148 1271 -1128 1275
rect -875 1271 -855 1275
rect -688 1271 -668 1275
rect -875 1263 -855 1267
rect -688 1263 -668 1267
rect -875 1255 -855 1259
rect -688 1255 -668 1259
rect -784 1249 -764 1253
rect -784 1241 -764 1245
rect -784 1233 -764 1237
rect -488 1198 -468 1202
rect -488 1190 -468 1194
rect -406 1192 -402 1212
rect -398 1192 -394 1212
rect -29 1199 -9 1203
rect -488 1182 -468 1186
rect -1476 1177 -1456 1181
rect -1149 1177 -1129 1181
rect -1476 1169 -1456 1173
rect -488 1174 -468 1178
rect -29 1191 -9 1195
rect -29 1183 -9 1187
rect -1149 1169 -1129 1173
rect -1582 1159 -1562 1163
rect -1476 1161 -1456 1165
rect -1255 1159 -1235 1163
rect -1582 1151 -1562 1155
rect -1149 1161 -1129 1165
rect -120 1165 -100 1169
rect 67 1165 87 1169
rect -120 1157 -100 1161
rect -1255 1151 -1235 1155
rect -1582 1143 -1562 1147
rect 67 1157 87 1161
rect -120 1149 -100 1153
rect 67 1149 87 1153
rect -1255 1143 -1235 1147
rect -29 1143 -9 1147
rect -1678 1111 -1674 1131
rect -1670 1111 -1666 1131
rect -1627 1111 -1623 1131
rect -1619 1111 -1615 1131
rect -1582 1112 -1562 1116
rect -1476 1112 -1456 1116
rect -1582 1104 -1562 1108
rect -1350 1111 -1346 1131
rect -1342 1111 -1338 1131
rect -1300 1111 -1296 1131
rect -1292 1111 -1288 1131
rect -408 1118 -404 1138
rect -400 1118 -396 1138
rect -29 1135 -9 1139
rect -29 1127 -9 1131
rect -1255 1112 -1235 1116
rect -1476 1104 -1456 1108
rect -1582 1096 -1562 1100
rect -1476 1096 -1456 1100
rect -1149 1112 -1129 1116
rect -1255 1104 -1235 1108
rect -481 1113 -461 1117
rect -1149 1104 -1129 1108
rect -1255 1096 -1235 1100
rect -481 1105 -461 1109
rect -1149 1096 -1129 1100
rect -481 1097 -461 1101
rect -292 1084 -232 1088
rect -292 1076 -232 1080
rect -190 1079 -186 1099
rect -182 1079 -178 1099
rect -292 1068 -232 1072
rect -292 1060 -232 1064
rect -891 1015 -871 1019
rect -891 1007 -871 1011
rect -1476 1002 -1456 1006
rect -1149 1002 -1129 1006
rect -1476 994 -1456 998
rect -797 1007 -793 1027
rect -789 1007 -785 1027
rect -891 999 -871 1003
rect -1149 994 -1129 998
rect -1582 984 -1562 988
rect -1476 986 -1456 990
rect -1255 984 -1235 988
rect -1582 976 -1562 980
rect -1149 986 -1129 990
rect -1255 976 -1235 980
rect -1582 968 -1562 972
rect -1255 968 -1235 972
rect -1678 936 -1674 956
rect -1670 936 -1666 956
rect -1627 936 -1623 956
rect -1619 936 -1615 956
rect -1582 937 -1562 941
rect -1476 937 -1456 941
rect -1582 929 -1562 933
rect -1350 936 -1346 956
rect -1342 936 -1338 956
rect -1300 936 -1296 956
rect -1292 936 -1288 956
rect -1255 937 -1235 941
rect -1476 929 -1456 933
rect -1582 921 -1562 925
rect -1476 921 -1456 925
rect -1149 937 -1129 941
rect -1255 929 -1235 933
rect -788 939 -768 943
rect -1149 929 -1129 933
rect -1255 921 -1235 925
rect -788 931 -768 935
rect -1149 921 -1129 925
rect -788 923 -768 927
rect -879 905 -859 909
rect -692 905 -672 909
rect -879 897 -859 901
rect -692 897 -672 901
rect -879 889 -859 893
rect -692 889 -672 893
rect -788 883 -768 887
rect 79 880 99 884
rect -788 875 -768 879
rect 79 872 99 876
rect -788 867 -768 871
rect 79 864 99 868
rect -448 848 -428 852
rect -448 840 -428 844
rect -356 839 -352 859
rect -348 839 -344 859
rect -227 847 -147 851
rect -227 839 -147 843
rect -448 832 -428 836
rect -1476 826 -1456 830
rect -1149 826 -1129 830
rect -1476 818 -1456 822
rect -448 824 -428 828
rect -1149 818 -1129 822
rect -1582 808 -1562 812
rect -1476 810 -1456 814
rect -104 836 -100 856
rect -96 836 -92 856
rect -12 846 8 850
rect 175 846 195 850
rect -12 838 8 842
rect -227 831 -147 835
rect -227 823 -147 827
rect -448 816 -428 820
rect -1255 808 -1235 812
rect -1582 800 -1562 804
rect -1149 810 -1129 814
rect 175 838 195 842
rect -12 830 8 834
rect 175 830 195 834
rect 79 824 99 828
rect -227 815 -147 819
rect 79 816 99 820
rect 79 808 99 812
rect -1255 800 -1235 804
rect -1582 792 -1562 796
rect -1255 792 -1235 796
rect -1678 760 -1674 780
rect -1670 760 -1666 780
rect -1627 760 -1623 780
rect -1619 760 -1615 780
rect -1582 761 -1562 765
rect -1476 761 -1456 765
rect -1582 753 -1562 757
rect -1350 760 -1346 780
rect -1342 760 -1338 780
rect -1300 760 -1296 780
rect -1292 760 -1288 780
rect -446 775 -426 779
rect -446 767 -426 771
rect -1255 761 -1235 765
rect -1476 753 -1456 757
rect -1582 745 -1562 749
rect -1476 745 -1456 749
rect -1149 761 -1129 765
rect -1255 753 -1235 757
rect -364 769 -360 789
rect -356 769 -352 789
rect -446 759 -426 763
rect -1149 753 -1129 757
rect -1255 745 -1235 749
rect -446 751 -426 755
rect -1149 745 -1129 749
rect -373 694 -369 714
rect -365 694 -361 714
rect -446 689 -426 693
rect -446 681 -426 685
rect -446 673 -426 677
rect -891 657 -871 661
rect -1476 651 -1456 655
rect -1149 651 -1129 655
rect -1476 643 -1456 647
rect -891 649 -871 653
rect -1149 643 -1129 647
rect -1582 633 -1562 637
rect -1476 635 -1456 639
rect -797 649 -793 669
rect -789 649 -785 669
rect -891 641 -871 645
rect -1255 633 -1235 637
rect -1582 625 -1562 629
rect -1149 635 -1129 639
rect -1255 625 -1235 629
rect -1582 617 -1562 621
rect -1255 617 -1235 621
rect -1678 585 -1674 605
rect -1670 585 -1666 605
rect -1627 585 -1623 605
rect -1619 585 -1615 605
rect -1582 586 -1562 590
rect -1476 586 -1456 590
rect -1582 578 -1562 582
rect -1350 585 -1346 605
rect -1342 585 -1338 605
rect -1300 585 -1296 605
rect -1292 585 -1288 605
rect -1255 586 -1235 590
rect -1476 578 -1456 582
rect -1582 570 -1562 574
rect -1476 570 -1456 574
rect -1149 586 -1129 590
rect -1255 578 -1235 582
rect -1149 578 -1129 582
rect -1255 570 -1235 574
rect -788 581 -768 585
rect -1149 570 -1129 574
rect -788 573 -768 577
rect -788 565 -768 569
rect -879 547 -859 551
rect -692 547 -672 551
rect -879 539 -859 543
rect -692 539 -672 543
rect -879 531 -859 535
rect -692 531 -672 535
rect -788 525 -768 529
rect -788 517 -768 521
rect -788 509 -768 513
rect -1475 345 -1455 349
rect -1148 345 -1128 349
rect -1475 337 -1455 341
rect -1148 337 -1128 341
rect -1581 327 -1561 331
rect -1475 329 -1455 333
rect -1254 327 -1234 331
rect -1581 319 -1561 323
rect -1148 329 -1128 333
rect -1254 319 -1234 323
rect -1581 311 -1561 315
rect -1254 311 -1234 315
rect -1677 279 -1673 299
rect -1669 279 -1665 299
rect -1626 279 -1622 299
rect -1618 279 -1614 299
rect -1581 280 -1561 284
rect -1475 280 -1455 284
rect -1581 272 -1561 276
rect -1349 279 -1345 299
rect -1341 279 -1337 299
rect -1299 279 -1295 299
rect -1291 279 -1287 299
rect -1254 280 -1234 284
rect -1475 272 -1455 276
rect -1581 264 -1561 268
rect -1475 264 -1455 268
rect -1148 280 -1128 284
rect -1254 272 -1234 276
rect -1148 272 -1128 276
rect -1254 264 -1234 268
rect -1148 264 -1128 268
rect -891 210 -871 214
rect -891 202 -871 206
rect -797 202 -793 222
rect -789 202 -785 222
rect -891 194 -871 198
rect -1476 170 -1456 174
rect -1149 170 -1129 174
rect -1476 162 -1456 166
rect -1149 162 -1129 166
rect -1582 152 -1562 156
rect -1476 154 -1456 158
rect -1255 152 -1235 156
rect -1582 144 -1562 148
rect -1149 154 -1129 158
rect -1255 144 -1235 148
rect -1582 136 -1562 140
rect -1255 136 -1235 140
rect -788 134 -768 138
rect -788 126 -768 130
rect -1678 104 -1674 124
rect -1670 104 -1666 124
rect -1627 104 -1623 124
rect -1619 104 -1615 124
rect -1582 105 -1562 109
rect -1476 105 -1456 109
rect -1582 97 -1562 101
rect -1350 104 -1346 124
rect -1342 104 -1338 124
rect -1300 104 -1296 124
rect -1292 104 -1288 124
rect -788 118 -768 122
rect -1255 105 -1235 109
rect -1476 97 -1456 101
rect -1582 89 -1562 93
rect -1476 89 -1456 93
rect -1149 105 -1129 109
rect -1255 97 -1235 101
rect -1149 97 -1129 101
rect -1255 89 -1235 93
rect -879 100 -859 104
rect -692 100 -672 104
rect -1149 89 -1129 93
rect -879 92 -859 96
rect -692 92 -672 96
rect -879 84 -859 88
rect -692 84 -672 88
rect -788 78 -768 82
rect -788 70 -768 74
rect -788 62 -768 66
rect -1476 -5 -1456 -1
rect -1149 -5 -1129 -1
rect -1476 -13 -1456 -9
rect -1149 -13 -1129 -9
rect -1582 -23 -1562 -19
rect -1476 -21 -1456 -17
rect -1255 -23 -1235 -19
rect -1582 -31 -1562 -27
rect -1149 -21 -1129 -17
rect -1255 -31 -1235 -27
rect -1582 -39 -1562 -35
rect -1255 -39 -1235 -35
rect -1678 -71 -1674 -51
rect -1670 -71 -1666 -51
rect -1627 -71 -1623 -51
rect -1619 -71 -1615 -51
rect -1582 -70 -1562 -66
rect -1476 -70 -1456 -66
rect -1582 -78 -1562 -74
rect -1350 -71 -1346 -51
rect -1342 -71 -1338 -51
rect -1300 -71 -1296 -51
rect -1292 -71 -1288 -51
rect -1255 -70 -1235 -66
rect -1476 -78 -1456 -74
rect -1582 -86 -1562 -82
rect -1476 -86 -1456 -82
rect -1149 -70 -1129 -66
rect -1255 -78 -1235 -74
rect -1149 -78 -1129 -74
rect -1255 -86 -1235 -82
rect -1149 -86 -1129 -82
rect -1476 -181 -1456 -177
rect -1149 -181 -1129 -177
rect -1476 -189 -1456 -185
rect -1149 -189 -1129 -185
rect -1582 -199 -1562 -195
rect -1476 -197 -1456 -193
rect -1255 -199 -1235 -195
rect -1582 -207 -1562 -203
rect -1149 -197 -1129 -193
rect -1255 -207 -1235 -203
rect -1582 -215 -1562 -211
rect -1255 -215 -1235 -211
rect -1678 -247 -1674 -227
rect -1670 -247 -1666 -227
rect -1627 -247 -1623 -227
rect -1619 -247 -1615 -227
rect -1582 -246 -1562 -242
rect -1476 -246 -1456 -242
rect -1582 -254 -1562 -250
rect -1350 -247 -1346 -227
rect -1342 -247 -1338 -227
rect -1300 -247 -1296 -227
rect -1292 -247 -1288 -227
rect -1255 -246 -1235 -242
rect -1476 -254 -1456 -250
rect -1582 -262 -1562 -258
rect -1476 -262 -1456 -258
rect -1149 -246 -1129 -242
rect -1255 -254 -1235 -250
rect -1149 -254 -1129 -250
rect -1255 -262 -1235 -258
rect -1149 -262 -1129 -258
rect -891 -293 -871 -289
rect -891 -301 -871 -297
rect -797 -301 -793 -281
rect -789 -301 -785 -281
rect -891 -309 -871 -305
rect -1476 -356 -1456 -352
rect -1149 -356 -1129 -352
rect -1476 -364 -1456 -360
rect -1149 -364 -1129 -360
rect -1582 -374 -1562 -370
rect -1476 -372 -1456 -368
rect -1255 -374 -1235 -370
rect -1582 -382 -1562 -378
rect -1149 -372 -1129 -368
rect -788 -369 -768 -365
rect -788 -377 -768 -373
rect -1255 -382 -1235 -378
rect -1582 -390 -1562 -386
rect -788 -385 -768 -381
rect -1255 -390 -1235 -386
rect -1678 -422 -1674 -402
rect -1670 -422 -1666 -402
rect -1627 -422 -1623 -402
rect -1619 -422 -1615 -402
rect -1582 -421 -1562 -417
rect -1476 -421 -1456 -417
rect -1582 -429 -1562 -425
rect -1350 -422 -1346 -402
rect -1342 -422 -1338 -402
rect -1300 -422 -1296 -402
rect -1292 -422 -1288 -402
rect -879 -403 -859 -399
rect -692 -403 -672 -399
rect -879 -411 -859 -407
rect -692 -411 -672 -407
rect -1255 -421 -1235 -417
rect -1476 -429 -1456 -425
rect -1582 -437 -1562 -433
rect -1476 -437 -1456 -433
rect -1149 -421 -1129 -417
rect -1255 -429 -1235 -425
rect -879 -419 -859 -415
rect -692 -419 -672 -415
rect -1149 -429 -1129 -425
rect -1255 -437 -1235 -433
rect -788 -425 -768 -421
rect -1149 -437 -1129 -433
rect -788 -433 -768 -429
rect -788 -441 -768 -437
<< polysilicon >>
rect -1487 1527 -1475 1529
rect -1455 1527 -1439 1529
rect -1419 1527 -1416 1529
rect -1160 1527 -1148 1529
rect -1128 1527 -1112 1529
rect -1092 1527 -1089 1529
rect -1487 1519 -1475 1521
rect -1455 1519 -1439 1521
rect -1419 1519 -1416 1521
rect -1160 1519 -1148 1521
rect -1128 1519 -1112 1521
rect -1092 1519 -1089 1521
rect -1593 1509 -1581 1511
rect -1561 1509 -1545 1511
rect -1525 1509 -1522 1511
rect -1266 1509 -1254 1511
rect -1234 1509 -1218 1511
rect -1198 1509 -1195 1511
rect -1593 1501 -1581 1503
rect -1561 1501 -1545 1503
rect -1525 1501 -1522 1503
rect -399 1508 -397 1511
rect -1266 1501 -1254 1503
rect -1234 1501 -1218 1503
rect -1198 1501 -1195 1503
rect -1672 1484 -1670 1487
rect -1621 1484 -1619 1487
rect -1344 1484 -1342 1487
rect -1294 1484 -1292 1487
rect -1672 1450 -1670 1464
rect -1621 1450 -1619 1464
rect -1593 1462 -1581 1464
rect -1561 1462 -1545 1464
rect -1525 1462 -1522 1464
rect -486 1480 -477 1482
rect -457 1480 -444 1482
rect -424 1480 -421 1482
rect -486 1472 -477 1474
rect -457 1472 -444 1474
rect -424 1472 -421 1474
rect -399 1472 -397 1488
rect -251 1473 -249 1476
rect -1487 1462 -1475 1464
rect -1455 1462 -1439 1464
rect -1419 1462 -1416 1464
rect -1593 1454 -1581 1456
rect -1561 1454 -1545 1456
rect -1525 1454 -1522 1456
rect -1487 1454 -1475 1456
rect -1455 1454 -1439 1456
rect -1419 1454 -1416 1456
rect -1344 1450 -1342 1464
rect -1294 1450 -1292 1464
rect -1266 1462 -1254 1464
rect -1234 1462 -1218 1464
rect -1198 1462 -1195 1464
rect -1160 1462 -1148 1464
rect -1128 1462 -1112 1464
rect -1092 1462 -1089 1464
rect -1266 1454 -1254 1456
rect -1234 1454 -1218 1456
rect -1198 1454 -1195 1456
rect -399 1459 -397 1462
rect -1160 1454 -1148 1456
rect -1128 1454 -1112 1456
rect -1092 1454 -1089 1456
rect -348 1444 -339 1446
rect -299 1444 -287 1446
rect -277 1444 -274 1446
rect -1672 1437 -1670 1440
rect -1621 1437 -1619 1440
rect -1344 1437 -1342 1440
rect -1294 1437 -1292 1440
rect -348 1436 -339 1438
rect -299 1436 -287 1438
rect -277 1436 -274 1438
rect -251 1437 -249 1453
rect -251 1424 -249 1427
rect -788 1393 -786 1396
rect -899 1378 -887 1380
rect -867 1378 -851 1380
rect -831 1378 -828 1380
rect -899 1370 -887 1372
rect -867 1370 -851 1372
rect -831 1370 -828 1372
rect -788 1359 -786 1373
rect -69 1363 -57 1365
rect -37 1363 -21 1365
rect -1 1363 2 1365
rect -1487 1349 -1475 1351
rect -1455 1349 -1439 1351
rect -1419 1349 -1416 1351
rect -1160 1349 -1148 1351
rect -1128 1349 -1112 1351
rect -1092 1349 -1089 1351
rect -69 1355 -57 1357
rect -37 1355 -21 1357
rect -1 1355 2 1357
rect -1487 1341 -1475 1343
rect -1455 1341 -1439 1343
rect -1419 1341 -1416 1343
rect -788 1346 -786 1349
rect -1160 1341 -1148 1343
rect -1128 1341 -1112 1343
rect -1092 1341 -1089 1343
rect -1593 1331 -1581 1333
rect -1561 1331 -1545 1333
rect -1525 1331 -1522 1333
rect -1266 1331 -1254 1333
rect -1234 1331 -1218 1333
rect -1198 1331 -1195 1333
rect -1593 1323 -1581 1325
rect -1561 1323 -1545 1325
rect -1525 1323 -1522 1325
rect -160 1329 -148 1331
rect -128 1329 -112 1331
rect -92 1329 -89 1331
rect -1266 1323 -1254 1325
rect -1234 1323 -1218 1325
rect -1198 1323 -1195 1325
rect 27 1329 39 1331
rect 59 1329 75 1331
rect 95 1329 98 1331
rect -160 1321 -148 1323
rect -128 1321 -112 1323
rect -92 1321 -89 1323
rect 27 1321 39 1323
rect 59 1321 75 1323
rect 95 1321 98 1323
rect -1672 1306 -1670 1309
rect -1621 1306 -1619 1309
rect -1344 1306 -1342 1309
rect -1294 1306 -1292 1309
rect -1672 1272 -1670 1286
rect -1621 1272 -1619 1286
rect -1593 1284 -1581 1286
rect -1561 1284 -1545 1286
rect -1525 1284 -1522 1286
rect -69 1307 -57 1309
rect -37 1307 -21 1309
rect -1 1307 2 1309
rect -796 1302 -784 1304
rect -764 1302 -748 1304
rect -728 1302 -725 1304
rect -69 1299 -57 1301
rect -37 1299 -21 1301
rect -1 1299 2 1301
rect -796 1294 -784 1296
rect -764 1294 -748 1296
rect -728 1294 -725 1296
rect -1487 1284 -1475 1286
rect -1455 1284 -1439 1286
rect -1419 1284 -1416 1286
rect -1593 1276 -1581 1278
rect -1561 1276 -1545 1278
rect -1525 1276 -1522 1278
rect -1487 1276 -1475 1278
rect -1455 1276 -1439 1278
rect -1419 1276 -1416 1278
rect -1344 1272 -1342 1286
rect -1294 1272 -1292 1286
rect -1266 1284 -1254 1286
rect -1234 1284 -1218 1286
rect -1198 1284 -1195 1286
rect -1160 1284 -1148 1286
rect -1128 1284 -1112 1286
rect -1092 1284 -1089 1286
rect -1266 1276 -1254 1278
rect -1234 1276 -1218 1278
rect -1198 1276 -1195 1278
rect -1160 1276 -1148 1278
rect -1128 1276 -1112 1278
rect -1092 1276 -1089 1278
rect -887 1268 -875 1270
rect -855 1268 -839 1270
rect -819 1268 -816 1270
rect -1672 1259 -1670 1262
rect -1621 1259 -1619 1262
rect -1344 1259 -1342 1262
rect -1294 1259 -1292 1262
rect -700 1268 -688 1270
rect -668 1268 -652 1270
rect -632 1268 -629 1270
rect -887 1260 -875 1262
rect -855 1260 -839 1262
rect -819 1260 -816 1262
rect -700 1260 -688 1262
rect -668 1260 -652 1262
rect -632 1260 -629 1262
rect -796 1246 -784 1248
rect -764 1246 -748 1248
rect -728 1246 -725 1248
rect -796 1238 -784 1240
rect -764 1238 -748 1240
rect -728 1238 -725 1240
rect -401 1212 -399 1215
rect -497 1195 -488 1197
rect -468 1195 -456 1197
rect -426 1195 -423 1197
rect -41 1196 -29 1198
rect -9 1196 7 1198
rect 27 1196 30 1198
rect -497 1187 -488 1189
rect -468 1187 -456 1189
rect -426 1187 -423 1189
rect -1488 1174 -1476 1176
rect -1456 1174 -1440 1176
rect -1420 1174 -1417 1176
rect -497 1179 -488 1181
rect -468 1179 -456 1181
rect -426 1179 -423 1181
rect -1161 1174 -1149 1176
rect -1129 1174 -1113 1176
rect -1093 1174 -1090 1176
rect -401 1176 -399 1192
rect -41 1188 -29 1190
rect -9 1188 7 1190
rect 27 1188 30 1190
rect -1488 1166 -1476 1168
rect -1456 1166 -1440 1168
rect -1420 1166 -1417 1168
rect -1161 1166 -1149 1168
rect -1129 1166 -1113 1168
rect -1093 1166 -1090 1168
rect -1594 1156 -1582 1158
rect -1562 1156 -1546 1158
rect -1526 1156 -1523 1158
rect -401 1163 -399 1166
rect -132 1162 -120 1164
rect -100 1162 -84 1164
rect -64 1162 -61 1164
rect -1267 1156 -1255 1158
rect -1235 1156 -1219 1158
rect -1199 1156 -1196 1158
rect -1594 1148 -1582 1150
rect -1562 1148 -1546 1150
rect -1526 1148 -1523 1150
rect 55 1162 67 1164
rect 87 1162 103 1164
rect 123 1162 126 1164
rect -132 1154 -120 1156
rect -100 1154 -84 1156
rect -64 1154 -61 1156
rect -1267 1148 -1255 1150
rect -1235 1148 -1219 1150
rect -1199 1148 -1196 1150
rect 55 1154 67 1156
rect 87 1154 103 1156
rect 123 1154 126 1156
rect -403 1138 -401 1141
rect -41 1140 -29 1142
rect -9 1140 7 1142
rect 27 1140 30 1142
rect -1673 1131 -1671 1134
rect -1622 1131 -1620 1134
rect -1345 1131 -1343 1134
rect -1295 1131 -1293 1134
rect -1673 1097 -1671 1111
rect -1622 1097 -1620 1111
rect -1594 1109 -1582 1111
rect -1562 1109 -1546 1111
rect -1526 1109 -1523 1111
rect -41 1132 -29 1134
rect -9 1132 7 1134
rect 27 1132 30 1134
rect -1488 1109 -1476 1111
rect -1456 1109 -1440 1111
rect -1420 1109 -1417 1111
rect -1594 1101 -1582 1103
rect -1562 1101 -1546 1103
rect -1526 1101 -1523 1103
rect -1488 1101 -1476 1103
rect -1456 1101 -1440 1103
rect -1420 1101 -1417 1103
rect -1345 1097 -1343 1111
rect -1295 1097 -1293 1111
rect -1267 1109 -1255 1111
rect -1235 1109 -1219 1111
rect -1199 1109 -1196 1111
rect -1161 1109 -1149 1111
rect -1129 1109 -1113 1111
rect -1093 1109 -1090 1111
rect -490 1110 -481 1112
rect -461 1110 -448 1112
rect -428 1110 -425 1112
rect -1267 1101 -1255 1103
rect -1235 1101 -1219 1103
rect -1199 1101 -1196 1103
rect -1161 1101 -1149 1103
rect -1129 1101 -1113 1103
rect -1093 1101 -1090 1103
rect -490 1102 -481 1104
rect -461 1102 -448 1104
rect -428 1102 -425 1104
rect -403 1102 -401 1118
rect -185 1099 -183 1102
rect -403 1089 -401 1092
rect -1673 1084 -1671 1087
rect -1622 1084 -1620 1087
rect -1345 1084 -1343 1087
rect -1295 1084 -1293 1087
rect -301 1081 -292 1083
rect -232 1081 -220 1083
rect -210 1081 -207 1083
rect -301 1073 -292 1075
rect -232 1073 -220 1075
rect -210 1073 -207 1075
rect -301 1065 -292 1067
rect -232 1065 -220 1067
rect -210 1065 -207 1067
rect -185 1063 -183 1079
rect -185 1050 -183 1053
rect -792 1027 -790 1030
rect -903 1012 -891 1014
rect -871 1012 -855 1014
rect -835 1012 -832 1014
rect -1488 999 -1476 1001
rect -1456 999 -1440 1001
rect -1420 999 -1417 1001
rect -903 1004 -891 1006
rect -871 1004 -855 1006
rect -835 1004 -832 1006
rect -1161 999 -1149 1001
rect -1129 999 -1113 1001
rect -1093 999 -1090 1001
rect -1488 991 -1476 993
rect -1456 991 -1440 993
rect -1420 991 -1417 993
rect -792 993 -790 1007
rect -1161 991 -1149 993
rect -1129 991 -1113 993
rect -1093 991 -1090 993
rect -1594 981 -1582 983
rect -1562 981 -1546 983
rect -1526 981 -1523 983
rect -1267 981 -1255 983
rect -1235 981 -1219 983
rect -1199 981 -1196 983
rect -1594 973 -1582 975
rect -1562 973 -1546 975
rect -1526 973 -1523 975
rect -792 980 -790 983
rect -1267 973 -1255 975
rect -1235 973 -1219 975
rect -1199 973 -1196 975
rect -1673 956 -1671 959
rect -1622 956 -1620 959
rect -1345 956 -1343 959
rect -1295 956 -1293 959
rect -1673 922 -1671 936
rect -1622 922 -1620 936
rect -1594 934 -1582 936
rect -1562 934 -1546 936
rect -1526 934 -1523 936
rect -1488 934 -1476 936
rect -1456 934 -1440 936
rect -1420 934 -1417 936
rect -1594 926 -1582 928
rect -1562 926 -1546 928
rect -1526 926 -1523 928
rect -1488 926 -1476 928
rect -1456 926 -1440 928
rect -1420 926 -1417 928
rect -1345 922 -1343 936
rect -1295 922 -1293 936
rect -1267 934 -1255 936
rect -1235 934 -1219 936
rect -1199 934 -1196 936
rect -1161 934 -1149 936
rect -1129 934 -1113 936
rect -1093 934 -1090 936
rect -800 936 -788 938
rect -768 936 -752 938
rect -732 936 -729 938
rect -1267 926 -1255 928
rect -1235 926 -1219 928
rect -1199 926 -1196 928
rect -1161 926 -1149 928
rect -1129 926 -1113 928
rect -1093 926 -1090 928
rect -800 928 -788 930
rect -768 928 -752 930
rect -732 928 -729 930
rect -1673 909 -1671 912
rect -1622 909 -1620 912
rect -1345 909 -1343 912
rect -1295 909 -1293 912
rect -891 902 -879 904
rect -859 902 -843 904
rect -823 902 -820 904
rect -704 902 -692 904
rect -672 902 -656 904
rect -636 902 -633 904
rect -891 894 -879 896
rect -859 894 -843 896
rect -823 894 -820 896
rect -704 894 -692 896
rect -672 894 -656 896
rect -636 894 -633 896
rect -800 880 -788 882
rect -768 880 -752 882
rect -732 880 -729 882
rect 67 877 79 879
rect 99 877 115 879
rect 135 877 138 879
rect -800 872 -788 874
rect -768 872 -752 874
rect -732 872 -729 874
rect 67 869 79 871
rect 99 869 115 871
rect 135 869 138 871
rect -351 859 -349 862
rect -457 845 -448 847
rect -428 845 -416 847
rect -376 845 -373 847
rect -99 856 -97 859
rect -236 844 -227 846
rect -147 844 -135 846
rect -125 844 -122 846
rect -457 837 -448 839
rect -428 837 -416 839
rect -376 837 -373 839
rect -1488 823 -1476 825
rect -1456 823 -1440 825
rect -1420 823 -1417 825
rect -457 829 -448 831
rect -428 829 -416 831
rect -376 829 -373 831
rect -1161 823 -1149 825
rect -1129 823 -1113 825
rect -1093 823 -1090 825
rect -1488 815 -1476 817
rect -1456 815 -1440 817
rect -1420 815 -1417 817
rect -351 823 -349 839
rect -236 836 -227 838
rect -147 836 -135 838
rect -125 836 -122 838
rect -24 843 -12 845
rect 8 843 24 845
rect 44 843 47 845
rect -236 828 -227 830
rect -147 828 -135 830
rect -125 828 -122 830
rect -457 821 -448 823
rect -428 821 -416 823
rect -376 821 -373 823
rect -1161 815 -1149 817
rect -1129 815 -1113 817
rect -1093 815 -1090 817
rect -1594 805 -1582 807
rect -1562 805 -1546 807
rect -1526 805 -1523 807
rect -236 820 -227 822
rect -147 820 -135 822
rect -125 820 -122 822
rect -99 820 -97 836
rect 163 843 175 845
rect 195 843 211 845
rect 231 843 234 845
rect -24 835 -12 837
rect 8 835 24 837
rect 44 835 47 837
rect 163 835 175 837
rect 195 835 211 837
rect 231 835 234 837
rect 67 821 79 823
rect 99 821 115 823
rect 135 821 138 823
rect -351 810 -349 813
rect 67 813 79 815
rect 99 813 115 815
rect 135 813 138 815
rect -99 807 -97 810
rect -1267 805 -1255 807
rect -1235 805 -1219 807
rect -1199 805 -1196 807
rect -1594 797 -1582 799
rect -1562 797 -1546 799
rect -1526 797 -1523 799
rect -1267 797 -1255 799
rect -1235 797 -1219 799
rect -1199 797 -1196 799
rect -359 789 -357 792
rect -1673 780 -1671 783
rect -1622 780 -1620 783
rect -1345 780 -1343 783
rect -1295 780 -1293 783
rect -1673 746 -1671 760
rect -1622 746 -1620 760
rect -1594 758 -1582 760
rect -1562 758 -1546 760
rect -1526 758 -1523 760
rect -455 772 -446 774
rect -426 772 -414 774
rect -384 772 -381 774
rect -1488 758 -1476 760
rect -1456 758 -1440 760
rect -1420 758 -1417 760
rect -1594 750 -1582 752
rect -1562 750 -1546 752
rect -1526 750 -1523 752
rect -1488 750 -1476 752
rect -1456 750 -1440 752
rect -1420 750 -1417 752
rect -1345 746 -1343 760
rect -1295 746 -1293 760
rect -1267 758 -1255 760
rect -1235 758 -1219 760
rect -1199 758 -1196 760
rect -455 764 -446 766
rect -426 764 -414 766
rect -384 764 -381 766
rect -1161 758 -1149 760
rect -1129 758 -1113 760
rect -1093 758 -1090 760
rect -1267 750 -1255 752
rect -1235 750 -1219 752
rect -1199 750 -1196 752
rect -455 756 -446 758
rect -426 756 -414 758
rect -384 756 -381 758
rect -1161 750 -1149 752
rect -1129 750 -1113 752
rect -1093 750 -1090 752
rect -359 753 -357 769
rect -359 740 -357 743
rect -1673 733 -1671 736
rect -1622 733 -1620 736
rect -1345 733 -1343 736
rect -1295 733 -1293 736
rect -368 714 -366 717
rect -455 686 -446 688
rect -426 686 -413 688
rect -393 686 -390 688
rect -455 678 -446 680
rect -426 678 -413 680
rect -393 678 -390 680
rect -368 678 -366 694
rect -792 669 -790 672
rect -1488 648 -1476 650
rect -1456 648 -1440 650
rect -1420 648 -1417 650
rect -903 654 -891 656
rect -871 654 -855 656
rect -835 654 -832 656
rect -1161 648 -1149 650
rect -1129 648 -1113 650
rect -1093 648 -1090 650
rect -1488 640 -1476 642
rect -1456 640 -1440 642
rect -1420 640 -1417 642
rect -368 665 -366 668
rect -903 646 -891 648
rect -871 646 -855 648
rect -835 646 -832 648
rect -1161 640 -1149 642
rect -1129 640 -1113 642
rect -1093 640 -1090 642
rect -1594 630 -1582 632
rect -1562 630 -1546 632
rect -1526 630 -1523 632
rect -792 635 -790 649
rect -1267 630 -1255 632
rect -1235 630 -1219 632
rect -1199 630 -1196 632
rect -1594 622 -1582 624
rect -1562 622 -1546 624
rect -1526 622 -1523 624
rect -1267 622 -1255 624
rect -1235 622 -1219 624
rect -1199 622 -1196 624
rect -792 622 -790 625
rect -1673 605 -1671 608
rect -1622 605 -1620 608
rect -1345 605 -1343 608
rect -1295 605 -1293 608
rect -1673 571 -1671 585
rect -1622 571 -1620 585
rect -1594 583 -1582 585
rect -1562 583 -1546 585
rect -1526 583 -1523 585
rect -1488 583 -1476 585
rect -1456 583 -1440 585
rect -1420 583 -1417 585
rect -1594 575 -1582 577
rect -1562 575 -1546 577
rect -1526 575 -1523 577
rect -1488 575 -1476 577
rect -1456 575 -1440 577
rect -1420 575 -1417 577
rect -1345 571 -1343 585
rect -1295 571 -1293 585
rect -1267 583 -1255 585
rect -1235 583 -1219 585
rect -1199 583 -1196 585
rect -1161 583 -1149 585
rect -1129 583 -1113 585
rect -1093 583 -1090 585
rect -1267 575 -1255 577
rect -1235 575 -1219 577
rect -1199 575 -1196 577
rect -800 578 -788 580
rect -768 578 -752 580
rect -732 578 -729 580
rect -1161 575 -1149 577
rect -1129 575 -1113 577
rect -1093 575 -1090 577
rect -800 570 -788 572
rect -768 570 -752 572
rect -732 570 -729 572
rect -1673 558 -1671 561
rect -1622 558 -1620 561
rect -1345 558 -1343 561
rect -1295 558 -1293 561
rect -891 544 -879 546
rect -859 544 -843 546
rect -823 544 -820 546
rect -704 544 -692 546
rect -672 544 -656 546
rect -636 544 -633 546
rect -891 536 -879 538
rect -859 536 -843 538
rect -823 536 -820 538
rect -704 536 -692 538
rect -672 536 -656 538
rect -636 536 -633 538
rect -800 522 -788 524
rect -768 522 -752 524
rect -732 522 -729 524
rect -800 514 -788 516
rect -768 514 -752 516
rect -732 514 -729 516
rect -1487 342 -1475 344
rect -1455 342 -1439 344
rect -1419 342 -1416 344
rect -1160 342 -1148 344
rect -1128 342 -1112 344
rect -1092 342 -1089 344
rect -1487 334 -1475 336
rect -1455 334 -1439 336
rect -1419 334 -1416 336
rect -1160 334 -1148 336
rect -1128 334 -1112 336
rect -1092 334 -1089 336
rect -1593 324 -1581 326
rect -1561 324 -1545 326
rect -1525 324 -1522 326
rect -1266 324 -1254 326
rect -1234 324 -1218 326
rect -1198 324 -1195 326
rect -1593 316 -1581 318
rect -1561 316 -1545 318
rect -1525 316 -1522 318
rect -1266 316 -1254 318
rect -1234 316 -1218 318
rect -1198 316 -1195 318
rect -1672 299 -1670 302
rect -1621 299 -1619 302
rect -1344 299 -1342 302
rect -1294 299 -1292 302
rect -1672 265 -1670 279
rect -1621 265 -1619 279
rect -1593 277 -1581 279
rect -1561 277 -1545 279
rect -1525 277 -1522 279
rect -1487 277 -1475 279
rect -1455 277 -1439 279
rect -1419 277 -1416 279
rect -1593 269 -1581 271
rect -1561 269 -1545 271
rect -1525 269 -1522 271
rect -1487 269 -1475 271
rect -1455 269 -1439 271
rect -1419 269 -1416 271
rect -1344 265 -1342 279
rect -1294 265 -1292 279
rect -1266 277 -1254 279
rect -1234 277 -1218 279
rect -1198 277 -1195 279
rect -1160 277 -1148 279
rect -1128 277 -1112 279
rect -1092 277 -1089 279
rect -1266 269 -1254 271
rect -1234 269 -1218 271
rect -1198 269 -1195 271
rect -1160 269 -1148 271
rect -1128 269 -1112 271
rect -1092 269 -1089 271
rect -1672 252 -1670 255
rect -1621 252 -1619 255
rect -1344 252 -1342 255
rect -1294 252 -1292 255
rect -792 222 -790 225
rect -903 207 -891 209
rect -871 207 -855 209
rect -835 207 -832 209
rect -903 199 -891 201
rect -871 199 -855 201
rect -835 199 -832 201
rect -792 188 -790 202
rect -792 175 -790 178
rect -1488 167 -1476 169
rect -1456 167 -1440 169
rect -1420 167 -1417 169
rect -1161 167 -1149 169
rect -1129 167 -1113 169
rect -1093 167 -1090 169
rect -1488 159 -1476 161
rect -1456 159 -1440 161
rect -1420 159 -1417 161
rect -1161 159 -1149 161
rect -1129 159 -1113 161
rect -1093 159 -1090 161
rect -1594 149 -1582 151
rect -1562 149 -1546 151
rect -1526 149 -1523 151
rect -1267 149 -1255 151
rect -1235 149 -1219 151
rect -1199 149 -1196 151
rect -1594 141 -1582 143
rect -1562 141 -1546 143
rect -1526 141 -1523 143
rect -1267 141 -1255 143
rect -1235 141 -1219 143
rect -1199 141 -1196 143
rect -800 131 -788 133
rect -768 131 -752 133
rect -732 131 -729 133
rect -1673 124 -1671 127
rect -1622 124 -1620 127
rect -1345 124 -1343 127
rect -1295 124 -1293 127
rect -1673 90 -1671 104
rect -1622 90 -1620 104
rect -1594 102 -1582 104
rect -1562 102 -1546 104
rect -1526 102 -1523 104
rect -800 123 -788 125
rect -768 123 -752 125
rect -732 123 -729 125
rect -1488 102 -1476 104
rect -1456 102 -1440 104
rect -1420 102 -1417 104
rect -1594 94 -1582 96
rect -1562 94 -1546 96
rect -1526 94 -1523 96
rect -1488 94 -1476 96
rect -1456 94 -1440 96
rect -1420 94 -1417 96
rect -1345 90 -1343 104
rect -1295 90 -1293 104
rect -1267 102 -1255 104
rect -1235 102 -1219 104
rect -1199 102 -1196 104
rect -1161 102 -1149 104
rect -1129 102 -1113 104
rect -1093 102 -1090 104
rect -1267 94 -1255 96
rect -1235 94 -1219 96
rect -1199 94 -1196 96
rect -891 97 -879 99
rect -859 97 -843 99
rect -823 97 -820 99
rect -1161 94 -1149 96
rect -1129 94 -1113 96
rect -1093 94 -1090 96
rect -704 97 -692 99
rect -672 97 -656 99
rect -636 97 -633 99
rect -891 89 -879 91
rect -859 89 -843 91
rect -823 89 -820 91
rect -704 89 -692 91
rect -672 89 -656 91
rect -636 89 -633 91
rect -1673 77 -1671 80
rect -1622 77 -1620 80
rect -1345 77 -1343 80
rect -1295 77 -1293 80
rect -800 75 -788 77
rect -768 75 -752 77
rect -732 75 -729 77
rect -800 67 -788 69
rect -768 67 -752 69
rect -732 67 -729 69
rect -1488 -8 -1476 -6
rect -1456 -8 -1440 -6
rect -1420 -8 -1417 -6
rect -1161 -8 -1149 -6
rect -1129 -8 -1113 -6
rect -1093 -8 -1090 -6
rect -1488 -16 -1476 -14
rect -1456 -16 -1440 -14
rect -1420 -16 -1417 -14
rect -1161 -16 -1149 -14
rect -1129 -16 -1113 -14
rect -1093 -16 -1090 -14
rect -1594 -26 -1582 -24
rect -1562 -26 -1546 -24
rect -1526 -26 -1523 -24
rect -1267 -26 -1255 -24
rect -1235 -26 -1219 -24
rect -1199 -26 -1196 -24
rect -1594 -34 -1582 -32
rect -1562 -34 -1546 -32
rect -1526 -34 -1523 -32
rect -1267 -34 -1255 -32
rect -1235 -34 -1219 -32
rect -1199 -34 -1196 -32
rect -1673 -51 -1671 -48
rect -1622 -51 -1620 -48
rect -1345 -51 -1343 -48
rect -1295 -51 -1293 -48
rect -1673 -85 -1671 -71
rect -1622 -85 -1620 -71
rect -1594 -73 -1582 -71
rect -1562 -73 -1546 -71
rect -1526 -73 -1523 -71
rect -1488 -73 -1476 -71
rect -1456 -73 -1440 -71
rect -1420 -73 -1417 -71
rect -1594 -81 -1582 -79
rect -1562 -81 -1546 -79
rect -1526 -81 -1523 -79
rect -1488 -81 -1476 -79
rect -1456 -81 -1440 -79
rect -1420 -81 -1417 -79
rect -1345 -85 -1343 -71
rect -1295 -85 -1293 -71
rect -1267 -73 -1255 -71
rect -1235 -73 -1219 -71
rect -1199 -73 -1196 -71
rect -1161 -73 -1149 -71
rect -1129 -73 -1113 -71
rect -1093 -73 -1090 -71
rect -1267 -81 -1255 -79
rect -1235 -81 -1219 -79
rect -1199 -81 -1196 -79
rect -1161 -81 -1149 -79
rect -1129 -81 -1113 -79
rect -1093 -81 -1090 -79
rect -1673 -98 -1671 -95
rect -1622 -98 -1620 -95
rect -1345 -98 -1343 -95
rect -1295 -98 -1293 -95
rect -1488 -184 -1476 -182
rect -1456 -184 -1440 -182
rect -1420 -184 -1417 -182
rect -1161 -184 -1149 -182
rect -1129 -184 -1113 -182
rect -1093 -184 -1090 -182
rect -1488 -192 -1476 -190
rect -1456 -192 -1440 -190
rect -1420 -192 -1417 -190
rect -1161 -192 -1149 -190
rect -1129 -192 -1113 -190
rect -1093 -192 -1090 -190
rect -1594 -202 -1582 -200
rect -1562 -202 -1546 -200
rect -1526 -202 -1523 -200
rect -1267 -202 -1255 -200
rect -1235 -202 -1219 -200
rect -1199 -202 -1196 -200
rect -1594 -210 -1582 -208
rect -1562 -210 -1546 -208
rect -1526 -210 -1523 -208
rect -1267 -210 -1255 -208
rect -1235 -210 -1219 -208
rect -1199 -210 -1196 -208
rect -1673 -227 -1671 -224
rect -1622 -227 -1620 -224
rect -1345 -227 -1343 -224
rect -1295 -227 -1293 -224
rect -1673 -261 -1671 -247
rect -1622 -261 -1620 -247
rect -1594 -249 -1582 -247
rect -1562 -249 -1546 -247
rect -1526 -249 -1523 -247
rect -1488 -249 -1476 -247
rect -1456 -249 -1440 -247
rect -1420 -249 -1417 -247
rect -1594 -257 -1582 -255
rect -1562 -257 -1546 -255
rect -1526 -257 -1523 -255
rect -1488 -257 -1476 -255
rect -1456 -257 -1440 -255
rect -1420 -257 -1417 -255
rect -1345 -261 -1343 -247
rect -1295 -261 -1293 -247
rect -1267 -249 -1255 -247
rect -1235 -249 -1219 -247
rect -1199 -249 -1196 -247
rect -1161 -249 -1149 -247
rect -1129 -249 -1113 -247
rect -1093 -249 -1090 -247
rect -1267 -257 -1255 -255
rect -1235 -257 -1219 -255
rect -1199 -257 -1196 -255
rect -1161 -257 -1149 -255
rect -1129 -257 -1113 -255
rect -1093 -257 -1090 -255
rect -1673 -274 -1671 -271
rect -1622 -274 -1620 -271
rect -1345 -274 -1343 -271
rect -1295 -274 -1293 -271
rect -792 -281 -790 -278
rect -903 -296 -891 -294
rect -871 -296 -855 -294
rect -835 -296 -832 -294
rect -903 -304 -891 -302
rect -871 -304 -855 -302
rect -835 -304 -832 -302
rect -792 -315 -790 -301
rect -792 -328 -790 -325
rect -1488 -359 -1476 -357
rect -1456 -359 -1440 -357
rect -1420 -359 -1417 -357
rect -1161 -359 -1149 -357
rect -1129 -359 -1113 -357
rect -1093 -359 -1090 -357
rect -1488 -367 -1476 -365
rect -1456 -367 -1440 -365
rect -1420 -367 -1417 -365
rect -1161 -367 -1149 -365
rect -1129 -367 -1113 -365
rect -1093 -367 -1090 -365
rect -1594 -377 -1582 -375
rect -1562 -377 -1546 -375
rect -1526 -377 -1523 -375
rect -800 -372 -788 -370
rect -768 -372 -752 -370
rect -732 -372 -729 -370
rect -1267 -377 -1255 -375
rect -1235 -377 -1219 -375
rect -1199 -377 -1196 -375
rect -1594 -385 -1582 -383
rect -1562 -385 -1546 -383
rect -1526 -385 -1523 -383
rect -800 -380 -788 -378
rect -768 -380 -752 -378
rect -732 -380 -729 -378
rect -1267 -385 -1255 -383
rect -1235 -385 -1219 -383
rect -1199 -385 -1196 -383
rect -1673 -402 -1671 -399
rect -1622 -402 -1620 -399
rect -1345 -402 -1343 -399
rect -1295 -402 -1293 -399
rect -1673 -436 -1671 -422
rect -1622 -436 -1620 -422
rect -1594 -424 -1582 -422
rect -1562 -424 -1546 -422
rect -1526 -424 -1523 -422
rect -891 -406 -879 -404
rect -859 -406 -843 -404
rect -823 -406 -820 -404
rect -704 -406 -692 -404
rect -672 -406 -656 -404
rect -636 -406 -633 -404
rect -891 -414 -879 -412
rect -859 -414 -843 -412
rect -823 -414 -820 -412
rect -1488 -424 -1476 -422
rect -1456 -424 -1440 -422
rect -1420 -424 -1417 -422
rect -1594 -432 -1582 -430
rect -1562 -432 -1546 -430
rect -1526 -432 -1523 -430
rect -1488 -432 -1476 -430
rect -1456 -432 -1440 -430
rect -1420 -432 -1417 -430
rect -1345 -436 -1343 -422
rect -1295 -436 -1293 -422
rect -1267 -424 -1255 -422
rect -1235 -424 -1219 -422
rect -1199 -424 -1196 -422
rect -704 -414 -692 -412
rect -672 -414 -656 -412
rect -636 -414 -633 -412
rect -1161 -424 -1149 -422
rect -1129 -424 -1113 -422
rect -1093 -424 -1090 -422
rect -1267 -432 -1255 -430
rect -1235 -432 -1219 -430
rect -1199 -432 -1196 -430
rect -800 -428 -788 -426
rect -768 -428 -752 -426
rect -732 -428 -729 -426
rect -1161 -432 -1149 -430
rect -1129 -432 -1113 -430
rect -1093 -432 -1090 -430
rect -800 -436 -788 -434
rect -768 -436 -752 -434
rect -732 -436 -729 -434
rect -1673 -449 -1671 -446
rect -1622 -449 -1620 -446
rect -1345 -449 -1343 -446
rect -1295 -449 -1293 -446
<< polycontact >>
rect -1491 1526 -1487 1530
rect -1491 1518 -1487 1522
rect -1164 1526 -1160 1530
rect -1597 1508 -1593 1512
rect -1164 1518 -1160 1522
rect -1597 1500 -1593 1504
rect -1270 1508 -1266 1512
rect -1270 1500 -1266 1504
rect -1676 1453 -1672 1457
rect -1625 1453 -1621 1457
rect -1597 1461 -1593 1465
rect -1597 1453 -1593 1457
rect -1491 1461 -1487 1465
rect -490 1479 -486 1483
rect -490 1471 -486 1475
rect -403 1475 -399 1479
rect -1491 1453 -1487 1457
rect -1348 1453 -1344 1457
rect -1298 1453 -1294 1457
rect -1270 1461 -1266 1465
rect -1270 1453 -1266 1457
rect -1164 1461 -1160 1465
rect -1164 1453 -1160 1457
rect -352 1443 -348 1447
rect -352 1435 -348 1439
rect -255 1440 -251 1444
rect -903 1377 -899 1381
rect -903 1369 -899 1373
rect -792 1362 -788 1366
rect -73 1362 -69 1366
rect -1491 1348 -1487 1352
rect -1491 1340 -1487 1344
rect -1164 1348 -1160 1352
rect -73 1354 -69 1358
rect -1597 1330 -1593 1334
rect -1164 1340 -1160 1344
rect -1597 1322 -1593 1326
rect -1270 1330 -1266 1334
rect -1270 1322 -1266 1326
rect -164 1328 -160 1332
rect -164 1320 -160 1324
rect 23 1328 27 1332
rect 23 1320 27 1324
rect -1676 1275 -1672 1279
rect -1625 1275 -1621 1279
rect -1597 1283 -1593 1287
rect -1597 1275 -1593 1279
rect -1491 1283 -1487 1287
rect -800 1301 -796 1305
rect -73 1306 -69 1310
rect -800 1293 -796 1297
rect -73 1298 -69 1302
rect -1491 1275 -1487 1279
rect -1348 1275 -1344 1279
rect -1298 1275 -1294 1279
rect -1270 1283 -1266 1287
rect -1270 1275 -1266 1279
rect -1164 1283 -1160 1287
rect -1164 1275 -1160 1279
rect -891 1267 -887 1271
rect -891 1259 -887 1263
rect -704 1267 -700 1271
rect -704 1259 -700 1263
rect -800 1245 -796 1249
rect -800 1237 -796 1241
rect -501 1194 -497 1198
rect -501 1186 -497 1190
rect -45 1195 -41 1199
rect -1492 1173 -1488 1177
rect -1492 1165 -1488 1169
rect -1165 1173 -1161 1177
rect -501 1178 -497 1182
rect -405 1179 -401 1183
rect -45 1187 -41 1191
rect -1598 1155 -1594 1159
rect -1165 1165 -1161 1169
rect -1598 1147 -1594 1151
rect -1271 1155 -1267 1159
rect -136 1161 -132 1165
rect -1271 1147 -1267 1151
rect -136 1153 -132 1157
rect 51 1161 55 1165
rect 51 1153 55 1157
rect -45 1139 -41 1143
rect -1677 1100 -1673 1104
rect -1626 1100 -1622 1104
rect -1598 1108 -1594 1112
rect -1598 1100 -1594 1104
rect -1492 1108 -1488 1112
rect -45 1131 -41 1135
rect -1492 1100 -1488 1104
rect -1349 1100 -1345 1104
rect -1299 1100 -1295 1104
rect -1271 1108 -1267 1112
rect -1271 1100 -1267 1104
rect -1165 1108 -1161 1112
rect -494 1109 -490 1113
rect -1165 1100 -1161 1104
rect -494 1101 -490 1105
rect -407 1105 -403 1109
rect -305 1080 -301 1084
rect -305 1072 -301 1076
rect -305 1064 -301 1068
rect -189 1066 -185 1070
rect -907 1011 -903 1015
rect -1492 998 -1488 1002
rect -1492 990 -1488 994
rect -1165 998 -1161 1002
rect -907 1003 -903 1007
rect -1598 980 -1594 984
rect -1165 990 -1161 994
rect -796 996 -792 1000
rect -1598 972 -1594 976
rect -1271 980 -1267 984
rect -1271 972 -1267 976
rect -1677 925 -1673 929
rect -1626 925 -1622 929
rect -1598 933 -1594 937
rect -1598 925 -1594 929
rect -1492 933 -1488 937
rect -1492 925 -1488 929
rect -1349 925 -1345 929
rect -1299 925 -1295 929
rect -1271 933 -1267 937
rect -1271 925 -1267 929
rect -1165 933 -1161 937
rect -804 935 -800 939
rect -1165 925 -1161 929
rect -804 927 -800 931
rect -895 901 -891 905
rect -895 893 -891 897
rect -708 901 -704 905
rect -708 893 -704 897
rect -804 879 -800 883
rect -804 871 -800 875
rect 63 876 67 880
rect 63 868 67 872
rect -461 844 -457 848
rect -461 836 -457 840
rect -240 843 -236 847
rect -1492 822 -1488 826
rect -1492 814 -1488 818
rect -1165 822 -1161 826
rect -461 828 -457 832
rect -1598 804 -1594 808
rect -1165 814 -1161 818
rect -461 820 -457 824
rect -355 826 -351 830
rect -240 835 -236 839
rect -28 842 -24 846
rect -240 827 -236 831
rect -1598 796 -1594 800
rect -1271 804 -1267 808
rect -240 819 -236 823
rect -103 823 -99 827
rect -28 834 -24 838
rect 159 842 163 846
rect 159 834 163 838
rect 63 820 67 824
rect 63 812 67 816
rect -1271 796 -1267 800
rect -1677 749 -1673 753
rect -1626 749 -1622 753
rect -1598 757 -1594 761
rect -1598 749 -1594 753
rect -1492 757 -1488 761
rect -459 771 -455 775
rect -1492 749 -1488 753
rect -1349 749 -1345 753
rect -1299 749 -1295 753
rect -1271 757 -1267 761
rect -1271 749 -1267 753
rect -1165 757 -1161 761
rect -459 763 -455 767
rect -1165 749 -1161 753
rect -459 755 -455 759
rect -363 756 -359 760
rect -459 685 -455 689
rect -459 677 -455 681
rect -372 681 -368 685
rect -1492 647 -1488 651
rect -1492 639 -1488 643
rect -1165 647 -1161 651
rect -907 653 -903 657
rect -1598 629 -1594 633
rect -1165 639 -1161 643
rect -907 645 -903 649
rect -1598 621 -1594 625
rect -1271 629 -1267 633
rect -796 638 -792 642
rect -1271 621 -1267 625
rect -1677 574 -1673 578
rect -1626 574 -1622 578
rect -1598 582 -1594 586
rect -1598 574 -1594 578
rect -1492 582 -1488 586
rect -1492 574 -1488 578
rect -1349 574 -1345 578
rect -1299 574 -1295 578
rect -1271 582 -1267 586
rect -1271 574 -1267 578
rect -1165 582 -1161 586
rect -1165 574 -1161 578
rect -804 577 -800 581
rect -804 569 -800 573
rect -895 543 -891 547
rect -895 535 -891 539
rect -708 543 -704 547
rect -708 535 -704 539
rect -804 521 -800 525
rect -804 513 -800 517
rect -1491 341 -1487 345
rect -1491 333 -1487 337
rect -1164 341 -1160 345
rect -1597 323 -1593 327
rect -1164 333 -1160 337
rect -1597 315 -1593 319
rect -1270 323 -1266 327
rect -1270 315 -1266 319
rect -1676 268 -1672 272
rect -1625 268 -1621 272
rect -1597 276 -1593 280
rect -1597 268 -1593 272
rect -1491 276 -1487 280
rect -1491 268 -1487 272
rect -1348 268 -1344 272
rect -1298 268 -1294 272
rect -1270 276 -1266 280
rect -1270 268 -1266 272
rect -1164 276 -1160 280
rect -1164 268 -1160 272
rect -907 206 -903 210
rect -907 198 -903 202
rect -796 191 -792 195
rect -1492 166 -1488 170
rect -1492 158 -1488 162
rect -1165 166 -1161 170
rect -1598 148 -1594 152
rect -1165 158 -1161 162
rect -1598 140 -1594 144
rect -1271 148 -1267 152
rect -1271 140 -1267 144
rect -804 130 -800 134
rect -1677 93 -1673 97
rect -1626 93 -1622 97
rect -1598 101 -1594 105
rect -1598 93 -1594 97
rect -1492 101 -1488 105
rect -804 122 -800 126
rect -1492 93 -1488 97
rect -1349 93 -1345 97
rect -1299 93 -1295 97
rect -1271 101 -1267 105
rect -1271 93 -1267 97
rect -1165 101 -1161 105
rect -1165 93 -1161 97
rect -895 96 -891 100
rect -895 88 -891 92
rect -708 96 -704 100
rect -708 88 -704 92
rect -804 74 -800 78
rect -804 66 -800 70
rect -1492 -9 -1488 -5
rect -1492 -17 -1488 -13
rect -1165 -9 -1161 -5
rect -1598 -27 -1594 -23
rect -1165 -17 -1161 -13
rect -1598 -35 -1594 -31
rect -1271 -27 -1267 -23
rect -1271 -35 -1267 -31
rect -1677 -82 -1673 -78
rect -1626 -82 -1622 -78
rect -1598 -74 -1594 -70
rect -1598 -82 -1594 -78
rect -1492 -74 -1488 -70
rect -1492 -82 -1488 -78
rect -1349 -82 -1345 -78
rect -1299 -82 -1295 -78
rect -1271 -74 -1267 -70
rect -1271 -82 -1267 -78
rect -1165 -74 -1161 -70
rect -1165 -82 -1161 -78
rect -1492 -185 -1488 -181
rect -1492 -193 -1488 -189
rect -1165 -185 -1161 -181
rect -1598 -203 -1594 -199
rect -1165 -193 -1161 -189
rect -1598 -211 -1594 -207
rect -1271 -203 -1267 -199
rect -1271 -211 -1267 -207
rect -1677 -258 -1673 -254
rect -1626 -258 -1622 -254
rect -1598 -250 -1594 -246
rect -1598 -258 -1594 -254
rect -1492 -250 -1488 -246
rect -1492 -258 -1488 -254
rect -1349 -258 -1345 -254
rect -1299 -258 -1295 -254
rect -1271 -250 -1267 -246
rect -1271 -258 -1267 -254
rect -1165 -250 -1161 -246
rect -1165 -258 -1161 -254
rect -907 -297 -903 -293
rect -907 -305 -903 -301
rect -796 -312 -792 -308
rect -1492 -360 -1488 -356
rect -1492 -368 -1488 -364
rect -1165 -360 -1161 -356
rect -1598 -378 -1594 -374
rect -1165 -368 -1161 -364
rect -1598 -386 -1594 -382
rect -1271 -378 -1267 -374
rect -804 -373 -800 -369
rect -1271 -386 -1267 -382
rect -804 -381 -800 -377
rect -1677 -433 -1673 -429
rect -1626 -433 -1622 -429
rect -1598 -425 -1594 -421
rect -1598 -433 -1594 -429
rect -1492 -425 -1488 -421
rect -895 -407 -891 -403
rect -895 -415 -891 -411
rect -708 -407 -704 -403
rect -1492 -433 -1488 -429
rect -1349 -433 -1345 -429
rect -1299 -433 -1295 -429
rect -1271 -425 -1267 -421
rect -1271 -433 -1267 -429
rect -1165 -425 -1161 -421
rect -708 -415 -704 -411
rect -1165 -433 -1161 -429
rect -804 -429 -800 -425
rect -804 -437 -800 -433
<< metal1 >>
rect -1533 1551 -1259 1554
rect -1533 1548 -1530 1551
rect -1263 1548 -1259 1551
rect -1703 1545 -1481 1548
rect -1751 1512 -1731 1521
rect -1590 1516 -1587 1545
rect -1484 1534 -1481 1545
rect -1263 1545 -1154 1548
rect -1447 1540 -1311 1544
rect -1484 1530 -1475 1534
rect -1553 1526 -1491 1530
rect -1590 1512 -1581 1516
rect -1751 1508 -1597 1512
rect -1751 1500 -1731 1508
rect -1683 1490 -1663 1494
rect -1677 1484 -1673 1490
rect -1669 1457 -1665 1464
rect -1652 1457 -1649 1499
rect -1737 1453 -1676 1457
rect -1669 1453 -1649 1457
rect -1642 1457 -1638 1508
rect -1627 1490 -1613 1494
rect -1626 1484 -1622 1490
rect -1618 1457 -1614 1464
rect -1601 1461 -1597 1504
rect -1590 1500 -1587 1512
rect -1553 1508 -1549 1526
rect -1519 1516 -1516 1522
rect -1525 1512 -1516 1516
rect -1561 1504 -1549 1508
rect -1553 1500 -1549 1504
rect -1590 1496 -1581 1500
rect -1553 1496 -1545 1500
rect -1590 1493 -1587 1496
rect -1519 1494 -1516 1512
rect -1484 1518 -1481 1530
rect -1447 1526 -1443 1540
rect -1419 1530 -1417 1534
rect -1455 1522 -1443 1526
rect -1447 1518 -1443 1522
rect -1491 1511 -1488 1518
rect -1484 1514 -1475 1518
rect -1447 1514 -1439 1518
rect -1484 1508 -1481 1514
rect -1409 1503 -1405 1540
rect -1491 1499 -1405 1503
rect -1553 1479 -1507 1483
rect -1590 1469 -1587 1472
rect -1590 1465 -1581 1469
rect -1642 1453 -1625 1457
rect -1618 1453 -1597 1457
rect -1590 1453 -1587 1465
rect -1553 1461 -1549 1479
rect -1519 1469 -1516 1471
rect -1525 1465 -1516 1469
rect -1561 1457 -1549 1461
rect -1553 1453 -1549 1457
rect -1771 1322 -1751 1343
rect -1771 1147 -1751 1168
rect -1771 972 -1751 993
rect -1771 796 -1751 817
rect -1771 621 -1751 642
rect -1771 315 -1751 336
rect -1771 140 -1751 161
rect -1771 -35 -1751 -14
rect -1771 -211 -1751 -190
rect -1771 -386 -1751 -365
rect -1737 -518 -1734 1453
rect -1669 1450 -1665 1453
rect -1618 1450 -1614 1453
rect -1590 1449 -1581 1453
rect -1553 1449 -1545 1453
rect -1590 1443 -1587 1449
rect -1677 1434 -1673 1440
rect -1626 1434 -1622 1440
rect -1519 1434 -1516 1465
rect -1511 1457 -1507 1479
rect -1491 1465 -1487 1499
rect -1484 1469 -1481 1475
rect -1484 1465 -1475 1469
rect -1511 1453 -1491 1457
rect -1484 1453 -1481 1465
rect -1447 1461 -1443 1491
rect -1399 1469 -1396 1530
rect -1315 1512 -1311 1540
rect -1263 1516 -1260 1545
rect -1157 1534 -1154 1545
rect -1120 1540 -212 1544
rect -1157 1530 -1148 1534
rect -1226 1526 -1164 1530
rect -1263 1512 -1254 1516
rect -1315 1508 -1270 1512
rect -1355 1490 -1331 1494
rect -1419 1465 -1396 1469
rect -1455 1457 -1443 1461
rect -1447 1453 -1443 1457
rect -1484 1449 -1475 1453
rect -1447 1449 -1439 1453
rect -1484 1443 -1481 1449
rect -1399 1434 -1396 1465
rect -1349 1484 -1345 1490
rect -1341 1457 -1337 1464
rect -1325 1457 -1320 1499
rect -1360 1453 -1348 1457
rect -1341 1453 -1320 1457
rect -1315 1457 -1311 1508
rect -1300 1490 -1286 1494
rect -1299 1484 -1295 1490
rect -1291 1457 -1287 1464
rect -1274 1461 -1270 1504
rect -1263 1500 -1260 1512
rect -1226 1508 -1222 1526
rect -1192 1516 -1189 1522
rect -1198 1512 -1189 1516
rect -1234 1504 -1222 1508
rect -1226 1500 -1222 1504
rect -1263 1496 -1254 1500
rect -1226 1496 -1218 1500
rect -1263 1493 -1260 1496
rect -1192 1494 -1189 1512
rect -1157 1518 -1154 1530
rect -1120 1526 -1116 1540
rect -1092 1530 -1090 1534
rect -1128 1522 -1116 1526
rect -1120 1518 -1116 1522
rect -1164 1511 -1161 1518
rect -1157 1514 -1148 1518
rect -1120 1514 -1112 1518
rect -1157 1508 -1154 1514
rect -1082 1503 -1078 1540
rect -1164 1499 -1078 1503
rect -1226 1479 -1180 1483
rect -1263 1469 -1260 1472
rect -1263 1465 -1254 1469
rect -1315 1453 -1298 1457
rect -1291 1453 -1270 1457
rect -1263 1453 -1260 1465
rect -1226 1461 -1222 1479
rect -1192 1469 -1189 1471
rect -1198 1465 -1189 1469
rect -1234 1457 -1222 1461
rect -1226 1453 -1222 1457
rect -1341 1450 -1337 1453
rect -1291 1450 -1287 1453
rect -1263 1449 -1254 1453
rect -1226 1449 -1218 1453
rect -1263 1443 -1260 1449
rect -1349 1434 -1345 1440
rect -1299 1434 -1295 1440
rect -1192 1434 -1189 1465
rect -1184 1457 -1180 1479
rect -1164 1465 -1160 1499
rect -1157 1469 -1154 1475
rect -1157 1465 -1148 1469
rect -1184 1453 -1164 1457
rect -1157 1453 -1154 1465
rect -1120 1461 -1116 1491
rect -1072 1469 -1069 1530
rect -1092 1465 -1069 1469
rect -1128 1457 -1116 1461
rect -1120 1453 -1116 1457
rect -1157 1449 -1148 1453
rect -1120 1449 -1112 1453
rect -1157 1443 -1154 1449
rect -1072 1434 -1069 1465
rect -567 1511 -525 1515
rect -1723 1431 -1069 1434
rect -1723 555 -1720 1431
rect -1708 1370 -1705 1412
rect -896 1399 -694 1403
rect -896 1385 -892 1399
rect -793 1393 -789 1399
rect -859 1388 -808 1392
rect -896 1381 -887 1385
rect -1070 1377 -903 1381
rect -1533 1373 -1259 1376
rect -1533 1370 -1530 1373
rect -1263 1370 -1259 1373
rect -1708 1367 -1481 1370
rect -1708 1195 -1705 1367
rect -1590 1338 -1587 1367
rect -1484 1356 -1481 1367
rect -1263 1367 -1154 1370
rect -1447 1362 -1311 1366
rect -1484 1352 -1475 1356
rect -1553 1348 -1491 1352
rect -1590 1334 -1581 1338
rect -1694 1330 -1597 1334
rect -1683 1312 -1663 1316
rect -1677 1306 -1673 1312
rect -1669 1279 -1665 1286
rect -1652 1279 -1649 1321
rect -1694 1275 -1676 1279
rect -1669 1275 -1649 1279
rect -1642 1279 -1638 1330
rect -1627 1312 -1613 1316
rect -1626 1306 -1622 1312
rect -1618 1279 -1614 1286
rect -1601 1283 -1597 1326
rect -1590 1322 -1587 1334
rect -1553 1330 -1549 1348
rect -1519 1338 -1516 1344
rect -1525 1334 -1516 1338
rect -1561 1326 -1549 1330
rect -1553 1322 -1549 1326
rect -1590 1318 -1581 1322
rect -1553 1318 -1545 1322
rect -1590 1315 -1587 1318
rect -1519 1316 -1516 1334
rect -1484 1340 -1481 1352
rect -1447 1348 -1443 1362
rect -1419 1352 -1417 1356
rect -1455 1344 -1443 1348
rect -1447 1340 -1443 1344
rect -1491 1333 -1488 1340
rect -1484 1336 -1475 1340
rect -1447 1336 -1439 1340
rect -1484 1330 -1481 1336
rect -1409 1325 -1405 1362
rect -1491 1321 -1405 1325
rect -1553 1301 -1507 1305
rect -1590 1291 -1587 1294
rect -1590 1287 -1581 1291
rect -1642 1275 -1625 1279
rect -1618 1275 -1597 1279
rect -1590 1275 -1587 1287
rect -1553 1283 -1549 1301
rect -1519 1291 -1516 1293
rect -1525 1287 -1516 1291
rect -1561 1279 -1549 1283
rect -1553 1275 -1549 1279
rect -1669 1272 -1665 1275
rect -1618 1272 -1614 1275
rect -1590 1271 -1581 1275
rect -1553 1271 -1545 1275
rect -1590 1265 -1587 1271
rect -1677 1256 -1673 1262
rect -1626 1256 -1622 1262
rect -1519 1256 -1516 1287
rect -1511 1279 -1507 1301
rect -1491 1287 -1487 1321
rect -1484 1291 -1481 1297
rect -1484 1287 -1475 1291
rect -1511 1275 -1491 1279
rect -1484 1275 -1481 1287
rect -1447 1283 -1443 1313
rect -1399 1291 -1396 1352
rect -1315 1334 -1311 1362
rect -1263 1338 -1260 1367
rect -1157 1356 -1154 1367
rect -1070 1366 -1066 1377
rect -1120 1362 -1066 1366
rect -1157 1352 -1148 1356
rect -1226 1348 -1164 1352
rect -1263 1334 -1254 1338
rect -1315 1330 -1270 1334
rect -1355 1312 -1331 1316
rect -1419 1287 -1396 1291
rect -1455 1279 -1443 1283
rect -1447 1275 -1443 1279
rect -1484 1271 -1475 1275
rect -1447 1271 -1439 1275
rect -1484 1265 -1481 1271
rect -1399 1256 -1396 1287
rect -1349 1306 -1345 1312
rect -1341 1279 -1337 1286
rect -1325 1279 -1320 1321
rect -1360 1275 -1348 1279
rect -1341 1275 -1320 1279
rect -1315 1279 -1311 1330
rect -1300 1312 -1286 1316
rect -1299 1306 -1295 1312
rect -1291 1279 -1287 1286
rect -1274 1283 -1270 1326
rect -1263 1322 -1260 1334
rect -1226 1330 -1222 1348
rect -1192 1338 -1189 1344
rect -1198 1334 -1189 1338
rect -1234 1326 -1222 1330
rect -1226 1322 -1222 1326
rect -1263 1318 -1254 1322
rect -1226 1318 -1218 1322
rect -1263 1315 -1260 1318
rect -1192 1316 -1189 1334
rect -1157 1340 -1154 1352
rect -1120 1348 -1116 1362
rect -1092 1352 -1090 1356
rect -1128 1344 -1116 1348
rect -1120 1340 -1116 1344
rect -1164 1333 -1161 1340
rect -1157 1336 -1148 1340
rect -1120 1336 -1112 1340
rect -1157 1330 -1154 1336
rect -1082 1325 -1078 1362
rect -1164 1321 -1078 1325
rect -1226 1301 -1180 1305
rect -1263 1291 -1260 1294
rect -1263 1287 -1254 1291
rect -1315 1275 -1298 1279
rect -1291 1275 -1270 1279
rect -1263 1275 -1260 1287
rect -1226 1283 -1222 1301
rect -1192 1291 -1189 1293
rect -1198 1287 -1189 1291
rect -1234 1279 -1222 1283
rect -1226 1275 -1222 1279
rect -1341 1272 -1337 1275
rect -1291 1272 -1287 1275
rect -1263 1271 -1254 1275
rect -1226 1271 -1218 1275
rect -1263 1265 -1260 1271
rect -1349 1256 -1345 1262
rect -1299 1256 -1295 1262
rect -1192 1256 -1189 1287
rect -1184 1279 -1180 1301
rect -1164 1287 -1160 1321
rect -1157 1291 -1154 1297
rect -1157 1287 -1148 1291
rect -1184 1275 -1164 1279
rect -1157 1275 -1154 1287
rect -1120 1283 -1116 1313
rect -1072 1291 -1069 1352
rect -1092 1287 -1069 1291
rect -1128 1279 -1116 1283
rect -1120 1275 -1116 1279
rect -1157 1271 -1148 1275
rect -1120 1271 -1112 1275
rect -1157 1265 -1154 1271
rect -1072 1256 -1069 1287
rect -1060 1273 -1056 1377
rect -1045 1369 -903 1373
rect -896 1369 -893 1381
rect -859 1377 -855 1388
rect -831 1381 -823 1385
rect -867 1373 -855 1377
rect -859 1369 -855 1373
rect -1677 1253 -1069 1256
rect -1045 1263 -1041 1369
rect -896 1365 -887 1369
rect -859 1365 -851 1369
rect -827 1347 -823 1381
rect -812 1366 -808 1388
rect -785 1366 -781 1373
rect -812 1362 -792 1366
rect -785 1362 -614 1366
rect -785 1359 -781 1362
rect -793 1347 -789 1349
rect -827 1343 -789 1347
rect -798 1339 -794 1343
rect -586 1339 -582 1455
rect -798 1335 -582 1339
rect -885 1323 -694 1327
rect -756 1312 -713 1316
rect -793 1305 -784 1309
rect -895 1301 -800 1305
rect -912 1273 -903 1277
rect -907 1271 -903 1273
rect -895 1271 -891 1301
rect -804 1282 -800 1297
rect -793 1293 -790 1305
rect -756 1301 -752 1312
rect -728 1305 -725 1309
rect -764 1297 -752 1301
rect -756 1293 -752 1297
rect -847 1278 -800 1282
rect -884 1271 -875 1275
rect -907 1267 -891 1271
rect -1045 1259 -891 1263
rect -884 1259 -881 1271
rect -847 1267 -843 1278
rect -819 1271 -815 1275
rect -855 1263 -843 1267
rect -847 1259 -843 1263
rect -1534 1198 -1260 1201
rect -1534 1195 -1531 1198
rect -1264 1195 -1260 1198
rect -1708 1192 -1482 1195
rect -1708 1020 -1705 1192
rect -1591 1163 -1588 1192
rect -1485 1181 -1482 1192
rect -1264 1192 -1155 1195
rect -1448 1187 -1312 1191
rect -1485 1177 -1476 1181
rect -1554 1173 -1492 1177
rect -1591 1159 -1582 1163
rect -1695 1155 -1598 1159
rect -1684 1137 -1664 1141
rect -1678 1131 -1674 1137
rect -1670 1104 -1666 1111
rect -1653 1104 -1650 1146
rect -1695 1100 -1677 1104
rect -1670 1100 -1650 1104
rect -1643 1104 -1639 1155
rect -1628 1137 -1614 1141
rect -1627 1131 -1623 1137
rect -1619 1104 -1615 1111
rect -1602 1108 -1598 1151
rect -1591 1147 -1588 1159
rect -1554 1155 -1550 1173
rect -1520 1163 -1517 1169
rect -1526 1159 -1517 1163
rect -1562 1151 -1550 1155
rect -1554 1147 -1550 1151
rect -1591 1143 -1582 1147
rect -1554 1143 -1546 1147
rect -1591 1140 -1588 1143
rect -1520 1141 -1517 1159
rect -1485 1165 -1482 1177
rect -1448 1173 -1444 1187
rect -1420 1177 -1418 1181
rect -1456 1169 -1444 1173
rect -1448 1165 -1444 1169
rect -1492 1158 -1489 1165
rect -1485 1161 -1476 1165
rect -1448 1161 -1440 1165
rect -1485 1155 -1482 1161
rect -1410 1150 -1406 1187
rect -1492 1146 -1406 1150
rect -1554 1126 -1508 1130
rect -1591 1116 -1588 1119
rect -1591 1112 -1582 1116
rect -1643 1100 -1626 1104
rect -1619 1100 -1598 1104
rect -1591 1100 -1588 1112
rect -1554 1108 -1550 1126
rect -1520 1116 -1517 1118
rect -1526 1112 -1517 1116
rect -1562 1104 -1550 1108
rect -1554 1100 -1550 1104
rect -1670 1097 -1666 1100
rect -1619 1097 -1615 1100
rect -1591 1096 -1582 1100
rect -1554 1096 -1546 1100
rect -1591 1090 -1588 1096
rect -1678 1081 -1674 1087
rect -1627 1081 -1623 1087
rect -1520 1081 -1517 1112
rect -1512 1104 -1508 1126
rect -1492 1112 -1488 1146
rect -1485 1116 -1482 1122
rect -1485 1112 -1476 1116
rect -1512 1100 -1492 1104
rect -1485 1100 -1482 1112
rect -1448 1108 -1444 1138
rect -1400 1116 -1397 1177
rect -1316 1159 -1312 1187
rect -1264 1163 -1261 1192
rect -1158 1181 -1155 1192
rect -1121 1187 -1061 1191
rect -1158 1177 -1149 1181
rect -1227 1173 -1165 1177
rect -1264 1159 -1255 1163
rect -1316 1155 -1271 1159
rect -1356 1137 -1332 1141
rect -1420 1112 -1397 1116
rect -1456 1104 -1444 1108
rect -1448 1100 -1444 1104
rect -1485 1096 -1476 1100
rect -1448 1096 -1440 1100
rect -1485 1090 -1482 1096
rect -1400 1081 -1397 1112
rect -1350 1131 -1346 1137
rect -1342 1104 -1338 1111
rect -1326 1104 -1321 1146
rect -1361 1100 -1349 1104
rect -1342 1100 -1321 1104
rect -1316 1104 -1312 1155
rect -1301 1137 -1287 1141
rect -1300 1131 -1296 1137
rect -1292 1104 -1288 1111
rect -1275 1108 -1271 1151
rect -1264 1147 -1261 1159
rect -1227 1155 -1223 1173
rect -1193 1163 -1190 1169
rect -1199 1159 -1190 1163
rect -1235 1151 -1223 1155
rect -1227 1147 -1223 1151
rect -1264 1143 -1255 1147
rect -1227 1143 -1219 1147
rect -1264 1140 -1261 1143
rect -1193 1141 -1190 1159
rect -1158 1165 -1155 1177
rect -1121 1173 -1117 1187
rect -1093 1177 -1091 1181
rect -1129 1169 -1117 1173
rect -1121 1165 -1117 1169
rect -1165 1158 -1162 1165
rect -1158 1161 -1149 1165
rect -1121 1161 -1113 1165
rect -1158 1155 -1155 1161
rect -1083 1150 -1079 1187
rect -1165 1146 -1079 1150
rect -1227 1126 -1181 1130
rect -1264 1116 -1261 1119
rect -1264 1112 -1255 1116
rect -1316 1100 -1299 1104
rect -1292 1100 -1271 1104
rect -1264 1100 -1261 1112
rect -1227 1108 -1223 1126
rect -1193 1116 -1190 1118
rect -1199 1112 -1190 1116
rect -1235 1104 -1223 1108
rect -1227 1100 -1223 1104
rect -1342 1097 -1338 1100
rect -1292 1097 -1288 1100
rect -1264 1096 -1255 1100
rect -1227 1096 -1219 1100
rect -1264 1090 -1261 1096
rect -1350 1081 -1346 1087
rect -1300 1081 -1296 1087
rect -1193 1081 -1190 1112
rect -1185 1104 -1181 1126
rect -1165 1112 -1161 1146
rect -1158 1116 -1155 1122
rect -1158 1112 -1149 1116
rect -1185 1100 -1165 1104
rect -1158 1100 -1155 1112
rect -1121 1108 -1117 1138
rect -1073 1116 -1070 1177
rect -1093 1112 -1070 1116
rect -1129 1104 -1117 1108
rect -1121 1100 -1117 1104
rect -1158 1096 -1149 1100
rect -1121 1096 -1113 1100
rect -1158 1090 -1155 1096
rect -1073 1081 -1070 1112
rect -1678 1078 -1070 1081
rect -1534 1023 -1260 1026
rect -1534 1020 -1531 1023
rect -1264 1020 -1260 1023
rect -1708 1017 -1482 1020
rect -1708 844 -1705 1017
rect -1591 988 -1588 1017
rect -1485 1006 -1482 1017
rect -1264 1017 -1155 1020
rect -1448 1012 -1312 1016
rect -1485 1002 -1476 1006
rect -1554 998 -1492 1002
rect -1591 984 -1582 988
rect -1695 980 -1598 984
rect -1684 962 -1664 966
rect -1678 956 -1674 962
rect -1670 929 -1666 936
rect -1653 929 -1650 971
rect -1695 925 -1677 929
rect -1670 925 -1650 929
rect -1643 929 -1639 980
rect -1628 962 -1614 966
rect -1627 956 -1623 962
rect -1619 929 -1615 936
rect -1602 933 -1598 976
rect -1591 972 -1588 984
rect -1554 980 -1550 998
rect -1520 988 -1517 994
rect -1526 984 -1517 988
rect -1562 976 -1550 980
rect -1554 972 -1550 976
rect -1591 968 -1582 972
rect -1554 968 -1546 972
rect -1591 965 -1588 968
rect -1520 966 -1517 984
rect -1485 990 -1482 1002
rect -1448 998 -1444 1012
rect -1420 1002 -1418 1006
rect -1456 994 -1444 998
rect -1448 990 -1444 994
rect -1492 983 -1489 990
rect -1485 986 -1476 990
rect -1448 986 -1440 990
rect -1485 980 -1482 986
rect -1410 975 -1406 1012
rect -1492 971 -1406 975
rect -1554 951 -1508 955
rect -1591 941 -1588 944
rect -1591 937 -1582 941
rect -1643 925 -1626 929
rect -1619 925 -1598 929
rect -1591 925 -1588 937
rect -1554 933 -1550 951
rect -1520 941 -1517 943
rect -1526 937 -1517 941
rect -1562 929 -1550 933
rect -1554 925 -1550 929
rect -1670 922 -1666 925
rect -1619 922 -1615 925
rect -1591 921 -1582 925
rect -1554 921 -1546 925
rect -1591 915 -1588 921
rect -1678 906 -1674 912
rect -1627 906 -1623 912
rect -1520 906 -1517 937
rect -1512 929 -1508 951
rect -1492 937 -1488 971
rect -1485 941 -1482 947
rect -1485 937 -1476 941
rect -1512 925 -1492 929
rect -1485 925 -1482 937
rect -1448 933 -1444 963
rect -1400 941 -1397 1002
rect -1316 984 -1312 1012
rect -1264 988 -1261 1017
rect -1158 1006 -1155 1017
rect -1121 1012 -1063 1016
rect -1158 1002 -1149 1006
rect -1227 998 -1165 1002
rect -1264 984 -1255 988
rect -1316 980 -1271 984
rect -1356 962 -1332 966
rect -1420 937 -1397 941
rect -1456 929 -1444 933
rect -1448 925 -1444 929
rect -1485 921 -1476 925
rect -1448 921 -1440 925
rect -1485 915 -1482 921
rect -1400 906 -1397 937
rect -1350 956 -1346 962
rect -1342 929 -1338 936
rect -1326 929 -1321 971
rect -1361 925 -1349 929
rect -1342 925 -1321 929
rect -1316 929 -1312 980
rect -1301 962 -1287 966
rect -1300 956 -1296 962
rect -1292 929 -1288 936
rect -1275 933 -1271 976
rect -1264 972 -1261 984
rect -1227 980 -1223 998
rect -1193 988 -1190 994
rect -1199 984 -1190 988
rect -1235 976 -1223 980
rect -1227 972 -1223 976
rect -1264 968 -1255 972
rect -1227 968 -1219 972
rect -1264 965 -1261 968
rect -1193 966 -1190 984
rect -1158 990 -1155 1002
rect -1121 998 -1117 1012
rect -1093 1002 -1091 1006
rect -1129 994 -1117 998
rect -1121 990 -1117 994
rect -1165 983 -1162 990
rect -1158 986 -1149 990
rect -1121 986 -1113 990
rect -1158 980 -1155 986
rect -1083 975 -1079 1012
rect -1165 971 -1079 975
rect -1227 951 -1181 955
rect -1264 941 -1261 944
rect -1264 937 -1255 941
rect -1316 925 -1299 929
rect -1292 925 -1271 929
rect -1264 925 -1261 937
rect -1227 933 -1223 951
rect -1193 941 -1190 943
rect -1199 937 -1190 941
rect -1235 929 -1223 933
rect -1227 925 -1223 929
rect -1342 922 -1338 925
rect -1292 922 -1288 925
rect -1264 921 -1255 925
rect -1227 921 -1219 925
rect -1264 915 -1261 921
rect -1350 906 -1346 912
rect -1300 906 -1296 912
rect -1193 906 -1190 937
rect -1185 929 -1181 951
rect -1165 937 -1161 971
rect -1158 941 -1155 947
rect -1158 937 -1149 941
rect -1185 925 -1165 929
rect -1158 925 -1155 937
rect -1121 933 -1117 963
rect -1073 941 -1070 1002
rect -1093 937 -1070 941
rect -1129 929 -1117 933
rect -1121 925 -1117 929
rect -1158 921 -1149 925
rect -1121 921 -1113 925
rect -1158 915 -1155 921
rect -1073 906 -1070 937
rect -1678 903 -1070 906
rect -1534 847 -1260 850
rect -1534 844 -1531 847
rect -1264 844 -1260 847
rect -1708 841 -1482 844
rect -1708 669 -1705 841
rect -1591 812 -1588 841
rect -1485 830 -1482 841
rect -1264 841 -1155 844
rect -1448 836 -1312 840
rect -1485 826 -1476 830
rect -1554 822 -1492 826
rect -1591 808 -1582 812
rect -1695 804 -1598 808
rect -1684 786 -1664 790
rect -1678 780 -1674 786
rect -1670 753 -1666 760
rect -1653 753 -1650 795
rect -1695 749 -1677 753
rect -1670 749 -1650 753
rect -1643 753 -1639 804
rect -1628 786 -1614 790
rect -1627 780 -1623 786
rect -1619 753 -1615 760
rect -1602 757 -1598 800
rect -1591 796 -1588 808
rect -1554 804 -1550 822
rect -1520 812 -1517 818
rect -1526 808 -1517 812
rect -1562 800 -1550 804
rect -1554 796 -1550 800
rect -1591 792 -1582 796
rect -1554 792 -1546 796
rect -1591 789 -1588 792
rect -1520 790 -1517 808
rect -1485 814 -1482 826
rect -1448 822 -1444 836
rect -1420 826 -1418 830
rect -1456 818 -1444 822
rect -1448 814 -1444 818
rect -1492 807 -1489 814
rect -1485 810 -1476 814
rect -1448 810 -1440 814
rect -1485 804 -1482 810
rect -1410 799 -1406 836
rect -1492 795 -1406 799
rect -1554 775 -1508 779
rect -1591 765 -1588 768
rect -1591 761 -1582 765
rect -1643 749 -1626 753
rect -1619 749 -1598 753
rect -1591 749 -1588 761
rect -1554 757 -1550 775
rect -1520 765 -1517 767
rect -1526 761 -1517 765
rect -1562 753 -1550 757
rect -1554 749 -1550 753
rect -1670 746 -1666 749
rect -1619 746 -1615 749
rect -1591 745 -1582 749
rect -1554 745 -1546 749
rect -1591 739 -1588 745
rect -1678 730 -1674 736
rect -1627 730 -1623 736
rect -1520 730 -1517 761
rect -1512 753 -1508 775
rect -1492 761 -1488 795
rect -1485 765 -1482 771
rect -1485 761 -1476 765
rect -1512 749 -1492 753
rect -1485 749 -1482 761
rect -1448 757 -1444 787
rect -1400 765 -1397 826
rect -1316 808 -1312 836
rect -1264 812 -1261 841
rect -1158 830 -1155 841
rect -1121 836 -1062 840
rect -1158 826 -1149 830
rect -1227 822 -1165 826
rect -1264 808 -1255 812
rect -1316 804 -1271 808
rect -1356 786 -1332 790
rect -1420 761 -1397 765
rect -1456 753 -1444 757
rect -1448 749 -1444 753
rect -1485 745 -1476 749
rect -1448 745 -1440 749
rect -1485 739 -1482 745
rect -1400 730 -1397 761
rect -1350 780 -1346 786
rect -1342 753 -1338 760
rect -1326 753 -1321 795
rect -1361 749 -1349 753
rect -1342 749 -1321 753
rect -1316 753 -1312 804
rect -1301 786 -1287 790
rect -1300 780 -1296 786
rect -1292 753 -1288 760
rect -1275 757 -1271 800
rect -1264 796 -1261 808
rect -1227 804 -1223 822
rect -1193 812 -1190 818
rect -1199 808 -1190 812
rect -1235 800 -1223 804
rect -1227 796 -1223 800
rect -1264 792 -1255 796
rect -1227 792 -1219 796
rect -1264 789 -1261 792
rect -1193 790 -1190 808
rect -1158 814 -1155 826
rect -1121 822 -1117 836
rect -1093 826 -1091 830
rect -1129 818 -1117 822
rect -1121 814 -1117 818
rect -1165 807 -1162 814
rect -1158 810 -1149 814
rect -1121 810 -1113 814
rect -1158 804 -1155 810
rect -1083 799 -1079 836
rect -1165 795 -1079 799
rect -1227 775 -1181 779
rect -1264 765 -1261 768
rect -1264 761 -1255 765
rect -1316 749 -1299 753
rect -1292 749 -1271 753
rect -1264 749 -1261 761
rect -1227 757 -1223 775
rect -1193 765 -1190 767
rect -1199 761 -1190 765
rect -1235 753 -1223 757
rect -1227 749 -1223 753
rect -1342 746 -1338 749
rect -1292 746 -1288 749
rect -1264 745 -1255 749
rect -1227 745 -1219 749
rect -1264 739 -1261 745
rect -1350 730 -1346 736
rect -1300 730 -1296 736
rect -1193 730 -1190 761
rect -1185 753 -1181 775
rect -1165 761 -1161 795
rect -1158 765 -1155 771
rect -1158 761 -1149 765
rect -1185 749 -1165 753
rect -1158 749 -1155 761
rect -1121 757 -1117 787
rect -1073 765 -1070 826
rect -1093 761 -1070 765
rect -1129 753 -1117 757
rect -1121 749 -1117 753
rect -1158 745 -1149 749
rect -1121 745 -1113 749
rect -1158 739 -1155 745
rect -1073 730 -1070 761
rect -1678 727 -1070 730
rect -1534 672 -1260 675
rect -1534 669 -1531 672
rect -1264 669 -1260 672
rect -1708 666 -1482 669
rect -1591 637 -1588 666
rect -1485 655 -1482 666
rect -1264 666 -1155 669
rect -1448 661 -1312 665
rect -1485 651 -1476 655
rect -1554 647 -1492 651
rect -1591 633 -1582 637
rect -1712 629 -1598 633
rect -1684 611 -1664 615
rect -1678 605 -1674 611
rect -1670 578 -1666 585
rect -1653 578 -1650 620
rect -1712 574 -1677 578
rect -1670 574 -1650 578
rect -1643 578 -1639 629
rect -1628 611 -1614 615
rect -1627 605 -1623 611
rect -1619 578 -1615 585
rect -1602 582 -1598 625
rect -1591 621 -1588 633
rect -1554 629 -1550 647
rect -1520 637 -1517 643
rect -1526 633 -1517 637
rect -1562 625 -1550 629
rect -1554 621 -1550 625
rect -1591 617 -1582 621
rect -1554 617 -1546 621
rect -1591 614 -1588 617
rect -1520 615 -1517 633
rect -1485 639 -1482 651
rect -1448 647 -1444 661
rect -1420 651 -1418 655
rect -1456 643 -1444 647
rect -1448 639 -1444 643
rect -1492 632 -1489 639
rect -1485 635 -1476 639
rect -1448 635 -1440 639
rect -1485 629 -1482 635
rect -1410 624 -1406 661
rect -1492 620 -1406 624
rect -1554 600 -1508 604
rect -1591 590 -1588 593
rect -1591 586 -1582 590
rect -1643 574 -1626 578
rect -1619 574 -1598 578
rect -1591 574 -1588 586
rect -1554 582 -1550 600
rect -1520 590 -1517 592
rect -1526 586 -1517 590
rect -1562 578 -1550 582
rect -1554 574 -1550 578
rect -1670 571 -1666 574
rect -1619 571 -1615 574
rect -1591 570 -1582 574
rect -1554 570 -1546 574
rect -1591 564 -1588 570
rect -1678 555 -1674 561
rect -1627 555 -1623 561
rect -1520 555 -1517 586
rect -1512 578 -1508 600
rect -1492 586 -1488 620
rect -1485 590 -1482 596
rect -1485 586 -1476 590
rect -1512 574 -1492 578
rect -1485 574 -1482 586
rect -1448 582 -1444 612
rect -1400 590 -1397 651
rect -1316 633 -1312 661
rect -1264 637 -1261 666
rect -1158 655 -1155 666
rect -1121 661 -1067 665
rect -1158 651 -1149 655
rect -1227 647 -1165 651
rect -1264 633 -1255 637
rect -1316 629 -1271 633
rect -1356 611 -1332 615
rect -1420 586 -1397 590
rect -1456 578 -1444 582
rect -1448 574 -1444 578
rect -1485 570 -1476 574
rect -1448 570 -1440 574
rect -1485 564 -1482 570
rect -1400 555 -1397 586
rect -1350 605 -1346 611
rect -1342 578 -1338 585
rect -1326 578 -1321 620
rect -1361 574 -1349 578
rect -1342 574 -1321 578
rect -1316 578 -1312 629
rect -1301 611 -1287 615
rect -1300 605 -1296 611
rect -1292 578 -1288 585
rect -1275 582 -1271 625
rect -1264 621 -1261 633
rect -1227 629 -1223 647
rect -1193 637 -1190 643
rect -1199 633 -1190 637
rect -1235 625 -1223 629
rect -1227 621 -1223 625
rect -1264 617 -1255 621
rect -1227 617 -1219 621
rect -1264 614 -1261 617
rect -1193 615 -1190 633
rect -1158 639 -1155 651
rect -1121 647 -1117 661
rect -1093 651 -1091 655
rect -1129 643 -1117 647
rect -1121 639 -1117 643
rect -1165 632 -1162 639
rect -1158 635 -1149 639
rect -1121 635 -1113 639
rect -1158 629 -1155 635
rect -1083 624 -1079 661
rect -1165 620 -1079 624
rect -1227 600 -1181 604
rect -1264 590 -1261 593
rect -1264 586 -1255 590
rect -1316 574 -1299 578
rect -1292 574 -1271 578
rect -1264 574 -1261 586
rect -1227 582 -1223 600
rect -1193 590 -1190 592
rect -1199 586 -1190 590
rect -1235 578 -1223 582
rect -1227 574 -1223 578
rect -1342 571 -1338 574
rect -1292 571 -1288 574
rect -1264 570 -1255 574
rect -1227 570 -1219 574
rect -1264 564 -1261 570
rect -1350 555 -1346 561
rect -1300 555 -1296 561
rect -1193 555 -1190 586
rect -1185 578 -1181 600
rect -1165 586 -1161 620
rect -1158 590 -1155 596
rect -1158 586 -1149 590
rect -1185 574 -1165 578
rect -1158 574 -1155 586
rect -1121 582 -1117 612
rect -1073 590 -1070 651
rect -1093 586 -1070 590
rect -1129 578 -1117 582
rect -1121 574 -1117 578
rect -1158 570 -1149 574
rect -1121 570 -1113 574
rect -1158 564 -1155 570
rect -1073 555 -1070 586
rect -1723 552 -1070 555
rect -1723 -452 -1720 552
rect -1708 363 -1705 507
rect -1533 366 -1259 369
rect -1533 363 -1530 366
rect -1263 363 -1259 366
rect -1708 360 -1481 363
rect -1708 188 -1705 360
rect -1590 331 -1587 360
rect -1484 349 -1481 360
rect -1263 360 -1154 363
rect -1447 355 -1311 359
rect -1484 345 -1475 349
rect -1553 341 -1491 345
rect -1590 327 -1581 331
rect -1694 323 -1597 327
rect -1683 305 -1663 309
rect -1677 299 -1673 305
rect -1669 272 -1665 279
rect -1652 272 -1649 314
rect -1694 268 -1676 272
rect -1669 268 -1649 272
rect -1642 272 -1638 323
rect -1627 305 -1613 309
rect -1626 299 -1622 305
rect -1618 272 -1614 279
rect -1601 276 -1597 319
rect -1590 315 -1587 327
rect -1553 323 -1549 341
rect -1519 331 -1516 337
rect -1525 327 -1516 331
rect -1561 319 -1549 323
rect -1553 315 -1549 319
rect -1590 311 -1581 315
rect -1553 311 -1545 315
rect -1590 308 -1587 311
rect -1519 309 -1516 327
rect -1484 333 -1481 345
rect -1447 341 -1443 355
rect -1419 345 -1417 349
rect -1455 337 -1443 341
rect -1447 333 -1443 337
rect -1491 326 -1488 333
rect -1484 329 -1475 333
rect -1447 329 -1439 333
rect -1484 323 -1481 329
rect -1409 318 -1405 355
rect -1491 314 -1405 318
rect -1553 294 -1507 298
rect -1590 284 -1587 287
rect -1590 280 -1581 284
rect -1642 268 -1625 272
rect -1618 268 -1597 272
rect -1590 268 -1587 280
rect -1553 276 -1549 294
rect -1519 284 -1516 286
rect -1525 280 -1516 284
rect -1561 272 -1549 276
rect -1553 268 -1549 272
rect -1669 265 -1665 268
rect -1618 265 -1614 268
rect -1590 264 -1581 268
rect -1553 264 -1545 268
rect -1590 258 -1587 264
rect -1677 249 -1673 255
rect -1626 249 -1622 255
rect -1519 249 -1516 280
rect -1511 272 -1507 294
rect -1491 280 -1487 314
rect -1484 284 -1481 290
rect -1484 280 -1475 284
rect -1511 268 -1491 272
rect -1484 268 -1481 280
rect -1447 276 -1443 306
rect -1399 284 -1396 345
rect -1315 327 -1311 355
rect -1263 331 -1260 360
rect -1157 349 -1154 360
rect -1045 359 -1041 1259
rect -895 1241 -891 1259
rect -884 1255 -875 1259
rect -847 1255 -839 1259
rect -804 1245 -800 1278
rect -793 1289 -784 1293
rect -756 1289 -748 1293
rect -793 1280 -789 1289
rect -793 1276 -744 1280
rect -793 1253 -789 1276
rect -717 1271 -713 1312
rect -698 1280 -694 1323
rect -660 1279 -614 1283
rect -697 1271 -688 1275
rect -717 1267 -704 1271
rect -717 1260 -704 1263
rect -756 1259 -704 1260
rect -697 1259 -694 1271
rect -660 1267 -656 1279
rect -632 1271 -628 1275
rect -668 1263 -656 1267
rect -660 1259 -656 1263
rect -756 1256 -713 1259
rect -793 1249 -784 1253
rect -895 1237 -800 1241
rect -793 1237 -790 1249
rect -756 1245 -752 1256
rect -697 1255 -688 1259
rect -660 1255 -652 1259
rect -728 1249 -718 1253
rect -764 1241 -752 1245
rect -756 1237 -752 1241
rect -793 1233 -784 1237
rect -756 1233 -748 1237
rect -722 1230 -718 1249
rect -628 1230 -624 1271
rect -586 1230 -582 1335
rect -790 1226 -582 1230
rect -916 1015 -911 1186
rect -900 1033 -698 1036
rect -900 1019 -896 1033
rect -797 1027 -793 1033
rect -863 1022 -812 1026
rect -900 1015 -891 1019
rect -916 1011 -907 1015
rect -1120 355 -1041 359
rect -1037 1003 -907 1007
rect -900 1003 -897 1015
rect -863 1011 -859 1022
rect -835 1015 -827 1019
rect -871 1007 -859 1011
rect -863 1003 -859 1007
rect -1037 897 -1033 1003
rect -900 999 -891 1003
rect -863 999 -855 1003
rect -831 981 -827 1015
rect -816 1000 -812 1022
rect -789 1000 -785 1007
rect -816 996 -796 1000
rect -789 996 -614 1000
rect -789 993 -785 996
rect -797 981 -793 983
rect -831 977 -793 981
rect -810 974 -806 977
rect -586 974 -582 1226
rect -810 970 -582 974
rect -889 957 -698 961
rect -760 946 -717 950
rect -797 939 -788 943
rect -899 935 -804 939
rect -899 905 -895 935
rect -808 916 -804 931
rect -797 927 -794 939
rect -760 935 -756 946
rect -732 939 -729 943
rect -768 931 -756 935
rect -760 927 -756 931
rect -851 912 -804 916
rect -888 905 -879 909
rect -928 904 -895 905
rect -933 901 -895 904
rect -1037 893 -895 897
rect -888 893 -885 905
rect -851 901 -847 912
rect -823 905 -819 909
rect -859 897 -847 901
rect -851 893 -847 897
rect -1157 345 -1148 349
rect -1226 341 -1164 345
rect -1263 327 -1254 331
rect -1315 323 -1270 327
rect -1355 305 -1331 309
rect -1419 280 -1396 284
rect -1455 272 -1443 276
rect -1447 268 -1443 272
rect -1484 264 -1475 268
rect -1447 264 -1439 268
rect -1484 258 -1481 264
rect -1399 249 -1396 280
rect -1349 299 -1345 305
rect -1341 272 -1337 279
rect -1325 272 -1320 314
rect -1360 268 -1348 272
rect -1341 268 -1320 272
rect -1315 272 -1311 323
rect -1300 305 -1286 309
rect -1299 299 -1295 305
rect -1291 272 -1287 279
rect -1274 276 -1270 319
rect -1263 315 -1260 327
rect -1226 323 -1222 341
rect -1192 331 -1189 337
rect -1198 327 -1189 331
rect -1234 319 -1222 323
rect -1226 315 -1222 319
rect -1263 311 -1254 315
rect -1226 311 -1218 315
rect -1263 308 -1260 311
rect -1192 309 -1189 327
rect -1157 333 -1154 345
rect -1120 341 -1116 355
rect -1092 345 -1090 349
rect -1128 337 -1116 341
rect -1120 333 -1116 337
rect -1164 326 -1161 333
rect -1157 329 -1148 333
rect -1120 329 -1112 333
rect -1157 323 -1154 329
rect -1082 318 -1078 355
rect -1164 314 -1078 318
rect -1226 294 -1180 298
rect -1263 284 -1260 287
rect -1263 280 -1254 284
rect -1315 268 -1298 272
rect -1291 268 -1270 272
rect -1263 268 -1260 280
rect -1226 276 -1222 294
rect -1192 284 -1189 286
rect -1198 280 -1189 284
rect -1234 272 -1222 276
rect -1226 268 -1222 272
rect -1341 265 -1337 268
rect -1291 265 -1287 268
rect -1263 264 -1254 268
rect -1226 264 -1218 268
rect -1263 258 -1260 264
rect -1349 249 -1345 255
rect -1299 249 -1295 255
rect -1192 249 -1189 280
rect -1184 272 -1180 294
rect -1164 280 -1160 314
rect -1157 284 -1154 290
rect -1157 280 -1148 284
rect -1184 268 -1164 272
rect -1157 268 -1154 280
rect -1120 276 -1116 306
rect -1072 284 -1069 345
rect -1092 280 -1069 284
rect -1128 272 -1116 276
rect -1120 268 -1116 272
rect -1157 264 -1148 268
rect -1120 264 -1112 268
rect -1157 258 -1154 264
rect -1072 249 -1069 280
rect -1677 246 -1069 249
rect -1534 191 -1260 194
rect -1534 188 -1531 191
rect -1264 188 -1260 191
rect -1708 185 -1482 188
rect -1708 13 -1705 185
rect -1591 156 -1588 185
rect -1485 174 -1482 185
rect -1264 185 -1155 188
rect -1448 180 -1312 184
rect -1485 170 -1476 174
rect -1554 166 -1492 170
rect -1591 152 -1582 156
rect -1695 148 -1598 152
rect -1684 130 -1664 134
rect -1678 124 -1674 130
rect -1670 97 -1666 104
rect -1653 97 -1650 139
rect -1695 93 -1677 97
rect -1670 93 -1650 97
rect -1643 97 -1639 148
rect -1628 130 -1614 134
rect -1627 124 -1623 130
rect -1619 97 -1615 104
rect -1602 101 -1598 144
rect -1591 140 -1588 152
rect -1554 148 -1550 166
rect -1520 156 -1517 162
rect -1526 152 -1517 156
rect -1562 144 -1550 148
rect -1554 140 -1550 144
rect -1591 136 -1582 140
rect -1554 136 -1546 140
rect -1591 133 -1588 136
rect -1520 134 -1517 152
rect -1485 158 -1482 170
rect -1448 166 -1444 180
rect -1420 170 -1418 174
rect -1456 162 -1444 166
rect -1448 158 -1444 162
rect -1492 151 -1489 158
rect -1485 154 -1476 158
rect -1448 154 -1440 158
rect -1485 148 -1482 154
rect -1410 143 -1406 180
rect -1492 139 -1406 143
rect -1554 119 -1508 123
rect -1591 109 -1588 112
rect -1591 105 -1582 109
rect -1643 93 -1626 97
rect -1619 93 -1598 97
rect -1591 93 -1588 105
rect -1554 101 -1550 119
rect -1520 109 -1517 111
rect -1526 105 -1517 109
rect -1562 97 -1550 101
rect -1554 93 -1550 97
rect -1670 90 -1666 93
rect -1619 90 -1615 93
rect -1591 89 -1582 93
rect -1554 89 -1546 93
rect -1591 83 -1588 89
rect -1678 74 -1674 80
rect -1627 74 -1623 80
rect -1520 74 -1517 105
rect -1512 97 -1508 119
rect -1492 105 -1488 139
rect -1485 109 -1482 115
rect -1485 105 -1476 109
rect -1512 93 -1492 97
rect -1485 93 -1482 105
rect -1448 101 -1444 131
rect -1400 109 -1397 170
rect -1316 152 -1312 180
rect -1264 156 -1261 185
rect -1158 174 -1155 185
rect -1037 184 -1033 893
rect -899 875 -895 893
rect -888 889 -879 893
rect -851 889 -843 893
rect -808 879 -804 912
rect -797 923 -788 927
rect -760 923 -752 927
rect -797 914 -793 923
rect -797 910 -748 914
rect -797 887 -793 910
rect -721 905 -717 946
rect -702 914 -698 957
rect -664 913 -614 917
rect -701 905 -692 909
rect -721 901 -708 905
rect -721 894 -708 897
rect -760 893 -708 894
rect -701 893 -698 905
rect -664 901 -660 913
rect -636 905 -632 909
rect -672 897 -660 901
rect -664 893 -660 897
rect -760 890 -717 893
rect -797 883 -788 887
rect -899 871 -804 875
rect -797 871 -794 883
rect -760 879 -756 890
rect -701 889 -692 893
rect -664 889 -656 893
rect -732 883 -722 887
rect -768 875 -756 879
rect -760 871 -756 875
rect -797 867 -788 871
rect -760 867 -752 871
rect -726 864 -722 883
rect -632 864 -628 905
rect -586 864 -582 970
rect -794 860 -582 864
rect -900 675 -698 678
rect -900 661 -896 675
rect -797 669 -793 675
rect -863 664 -812 668
rect -900 657 -891 661
rect -944 653 -907 657
rect -1121 180 -1033 184
rect -1019 645 -907 649
rect -900 645 -897 657
rect -863 653 -859 664
rect -835 657 -827 661
rect -871 649 -859 653
rect -863 645 -859 649
rect -1019 539 -1015 645
rect -900 641 -891 645
rect -863 641 -855 645
rect -831 623 -827 657
rect -816 642 -812 664
rect -789 642 -785 649
rect -816 638 -796 642
rect -789 638 -614 642
rect -789 635 -785 638
rect -797 623 -793 625
rect -831 619 -793 623
rect -808 615 -804 619
rect -586 615 -582 860
rect -567 865 -563 1511
rect -515 1483 -511 1540
rect -494 1511 -353 1514
rect -483 1487 -480 1511
rect -404 1508 -400 1511
rect -451 1490 -411 1494
rect -451 1487 -447 1490
rect -483 1483 -477 1487
rect -451 1483 -444 1487
rect -515 1479 -490 1483
rect -515 1471 -490 1475
rect -483 1471 -480 1483
rect -451 1479 -447 1483
rect -415 1479 -411 1490
rect -396 1479 -392 1488
rect -356 1479 -353 1511
rect -457 1475 -447 1479
rect -415 1475 -403 1479
rect -396 1475 -367 1479
rect -356 1476 -223 1479
rect -396 1472 -392 1475
rect -548 1354 -528 1375
rect -548 1284 -528 1292
rect -515 1284 -511 1471
rect -483 1467 -477 1471
rect -424 1467 -418 1471
rect -421 1459 -418 1467
rect -404 1459 -400 1462
rect -494 1456 -377 1459
rect -380 1425 -377 1456
rect -371 1447 -367 1475
rect -371 1443 -352 1447
rect -371 1435 -352 1439
rect -345 1435 -342 1476
rect -256 1473 -252 1476
rect -293 1454 -265 1457
rect -293 1451 -290 1454
rect -299 1447 -290 1451
rect -293 1443 -290 1447
rect -293 1439 -287 1443
rect -274 1435 -271 1451
rect -268 1444 -265 1454
rect -248 1444 -244 1453
rect -268 1440 -255 1444
rect -248 1440 -241 1444
rect -248 1437 -244 1440
rect -371 1366 -368 1435
rect -345 1431 -339 1435
rect -277 1431 -271 1435
rect -274 1424 -271 1431
rect -256 1424 -252 1427
rect -356 1421 -236 1424
rect -497 1363 -321 1366
rect -324 1292 -321 1363
rect -239 1293 -236 1421
rect -226 1388 -223 1476
rect -216 1332 -212 1540
rect -196 1384 33 1388
rect -29 1373 14 1377
rect -66 1366 -57 1370
rect -168 1362 -73 1366
rect -168 1332 -164 1362
rect -77 1343 -73 1358
rect -66 1354 -63 1366
rect -29 1362 -25 1373
rect -1 1366 2 1370
rect -37 1358 -25 1362
rect -29 1354 -25 1358
rect -120 1339 -73 1343
rect -157 1332 -148 1336
rect -216 1328 -164 1332
rect -191 1320 -164 1324
rect -157 1320 -154 1332
rect -120 1328 -116 1339
rect -92 1332 -88 1336
rect -128 1324 -116 1328
rect -120 1320 -116 1324
rect -239 1290 -206 1293
rect -191 1284 -187 1320
rect -168 1302 -164 1320
rect -157 1316 -148 1320
rect -120 1316 -112 1320
rect -77 1306 -73 1339
rect -66 1350 -57 1354
rect -29 1350 -21 1354
rect -66 1341 -62 1350
rect -66 1337 -17 1341
rect -66 1314 -62 1337
rect 10 1332 14 1373
rect 29 1341 33 1384
rect 117 1344 137 1353
rect 67 1340 137 1344
rect 30 1332 39 1336
rect 10 1328 23 1332
rect 10 1321 23 1324
rect -29 1320 23 1321
rect 30 1320 33 1332
rect 67 1328 71 1340
rect 95 1332 99 1336
rect 117 1332 137 1340
rect 59 1324 71 1328
rect 67 1320 71 1324
rect -29 1317 14 1320
rect -66 1310 -57 1314
rect -168 1298 -73 1302
rect -66 1298 -63 1310
rect -29 1306 -25 1317
rect 30 1316 39 1320
rect 67 1316 75 1320
rect -1 1310 9 1314
rect -37 1302 -25 1306
rect -29 1298 -25 1302
rect -66 1294 -57 1298
rect -29 1294 -21 1298
rect 5 1291 9 1310
rect 99 1291 103 1332
rect -175 1288 103 1291
rect -548 1280 -187 1284
rect -548 1271 -528 1280
rect -515 1266 -511 1280
rect -534 1262 -511 1266
rect -534 1190 -530 1262
rect -265 1258 -262 1268
rect -520 1255 -262 1258
rect -520 1198 -517 1255
rect -502 1215 -334 1218
rect -520 1194 -501 1198
rect -494 1194 -491 1215
rect -406 1212 -402 1215
rect -462 1205 -412 1208
rect -462 1202 -459 1205
rect -468 1198 -456 1202
rect -494 1190 -488 1194
rect -534 1186 -501 1190
rect -513 1178 -501 1182
rect -494 1178 -491 1190
rect -463 1186 -459 1198
rect -468 1182 -459 1186
rect -423 1178 -420 1202
rect -415 1183 -412 1205
rect -398 1183 -394 1192
rect -415 1179 -405 1183
rect -398 1179 -338 1183
rect -513 1105 -510 1178
rect -494 1174 -488 1178
rect -426 1174 -420 1178
rect -398 1176 -394 1179
rect -423 1163 -420 1174
rect -406 1163 -402 1166
rect -342 1163 -338 1179
rect -500 1160 -394 1163
rect -324 1155 -321 1243
rect -309 1217 61 1221
rect -506 1152 -321 1155
rect -506 1113 -503 1152
rect -309 1144 -306 1217
rect -1 1206 42 1210
rect -38 1199 -29 1203
rect -140 1195 -45 1199
rect -241 1165 -236 1167
rect -140 1165 -136 1195
rect -49 1176 -45 1191
rect -38 1187 -35 1199
rect -1 1195 3 1206
rect 27 1199 30 1203
rect -9 1191 3 1195
rect -1 1187 3 1191
rect -92 1172 -45 1176
rect -129 1165 -120 1169
rect -241 1161 -136 1165
rect -487 1141 -306 1144
rect -487 1117 -484 1141
rect -408 1138 -404 1141
rect -455 1120 -415 1124
rect -455 1117 -451 1120
rect -487 1113 -481 1117
rect -455 1113 -448 1117
rect -506 1109 -494 1113
rect -513 1101 -494 1105
rect -487 1101 -484 1113
rect -455 1109 -451 1113
rect -419 1109 -415 1120
rect -341 1126 -338 1133
rect -341 1123 -327 1126
rect -400 1109 -396 1118
rect -461 1105 -451 1109
rect -419 1105 -407 1109
rect -400 1105 -343 1109
rect -400 1102 -396 1105
rect -548 989 -528 1010
rect -548 917 -528 926
rect -513 917 -510 1101
rect -487 1097 -481 1101
rect -428 1097 -422 1101
rect -425 1089 -422 1097
rect -408 1089 -404 1092
rect -425 1086 -404 1089
rect -347 1076 -343 1105
rect -330 1084 -327 1123
rect -309 1105 -306 1141
rect -140 1135 -136 1157
rect -129 1153 -126 1165
rect -92 1161 -88 1172
rect -64 1165 -60 1169
rect -100 1157 -88 1161
rect -92 1153 -88 1157
rect -129 1149 -120 1153
rect -92 1149 -84 1153
rect -49 1139 -45 1172
rect -38 1183 -29 1187
rect -1 1183 7 1187
rect -38 1174 -34 1183
rect -38 1170 11 1174
rect -38 1147 -34 1170
rect 38 1165 42 1206
rect 57 1174 61 1217
rect 141 1177 161 1186
rect 95 1173 161 1177
rect 58 1165 67 1169
rect 38 1161 51 1165
rect 38 1154 51 1157
rect -1 1153 51 1154
rect 58 1153 61 1165
rect 95 1161 99 1173
rect 123 1165 127 1169
rect 141 1165 161 1173
rect 87 1157 99 1161
rect 95 1153 99 1157
rect -1 1150 42 1153
rect -38 1143 -29 1147
rect -140 1131 -45 1135
rect -38 1131 -35 1143
rect -1 1139 3 1150
rect 58 1149 67 1153
rect 95 1149 103 1153
rect 27 1143 37 1147
rect -9 1135 3 1139
rect -1 1131 3 1135
rect -38 1127 -29 1131
rect -1 1127 7 1131
rect 33 1124 37 1143
rect 127 1124 131 1165
rect -148 1120 131 1124
rect -309 1102 -172 1105
rect -330 1080 -305 1084
rect -347 1072 -305 1076
rect -467 1064 -305 1068
rect -298 1064 -295 1102
rect -190 1099 -186 1102
rect -226 1091 -196 1094
rect -226 1088 -223 1091
rect -232 1084 -220 1088
rect -226 1072 -223 1084
rect -207 1080 -204 1088
rect -210 1076 -204 1080
rect -226 1068 -220 1072
rect -207 1064 -204 1076
rect -199 1070 -196 1091
rect -182 1070 -178 1079
rect -199 1066 -189 1070
rect -182 1066 -60 1070
rect -467 1001 -463 1064
rect -420 1031 -416 1064
rect -298 1060 -292 1064
rect -210 1060 -204 1064
rect -182 1063 -178 1066
rect -298 1054 -295 1060
rect -207 1050 -204 1060
rect -190 1050 -186 1053
rect -357 1047 -178 1050
rect -420 1027 -180 1031
rect -175 1027 -137 1030
rect -490 986 -159 989
rect -490 917 -487 986
rect -140 950 -137 1027
rect -548 914 -487 917
rect -305 947 -137 950
rect -548 905 -528 914
rect -567 862 -320 865
rect -808 611 -582 615
rect -889 599 -698 603
rect -760 588 -717 592
rect -797 581 -788 585
rect -899 577 -804 581
rect -899 547 -895 577
rect -808 558 -804 573
rect -797 569 -794 581
rect -760 577 -756 588
rect -732 581 -729 585
rect -768 573 -756 577
rect -760 569 -756 573
rect -851 554 -804 558
rect -888 547 -879 551
rect -944 543 -895 547
rect -1019 535 -895 539
rect -888 535 -885 547
rect -851 543 -847 554
rect -823 547 -819 551
rect -859 539 -847 543
rect -851 535 -847 539
rect -1158 170 -1149 174
rect -1227 166 -1165 170
rect -1264 152 -1255 156
rect -1316 148 -1271 152
rect -1356 130 -1332 134
rect -1420 105 -1397 109
rect -1456 97 -1444 101
rect -1448 93 -1444 97
rect -1485 89 -1476 93
rect -1448 89 -1440 93
rect -1485 83 -1482 89
rect -1400 74 -1397 105
rect -1350 124 -1346 130
rect -1342 97 -1338 104
rect -1326 97 -1321 139
rect -1361 93 -1349 97
rect -1342 93 -1321 97
rect -1316 97 -1312 148
rect -1301 130 -1287 134
rect -1300 124 -1296 130
rect -1292 97 -1288 104
rect -1275 101 -1271 144
rect -1264 140 -1261 152
rect -1227 148 -1223 166
rect -1193 156 -1190 162
rect -1199 152 -1190 156
rect -1235 144 -1223 148
rect -1227 140 -1223 144
rect -1264 136 -1255 140
rect -1227 136 -1219 140
rect -1264 133 -1261 136
rect -1193 134 -1190 152
rect -1158 158 -1155 170
rect -1121 166 -1117 180
rect -1093 170 -1091 174
rect -1129 162 -1117 166
rect -1121 158 -1117 162
rect -1165 151 -1162 158
rect -1158 154 -1149 158
rect -1121 154 -1113 158
rect -1158 148 -1155 154
rect -1083 143 -1079 180
rect -1165 139 -1079 143
rect -1227 119 -1181 123
rect -1264 109 -1261 112
rect -1264 105 -1255 109
rect -1316 93 -1299 97
rect -1292 93 -1271 97
rect -1264 93 -1261 105
rect -1227 101 -1223 119
rect -1193 109 -1190 111
rect -1199 105 -1190 109
rect -1235 97 -1223 101
rect -1227 93 -1223 97
rect -1342 90 -1338 93
rect -1292 90 -1288 93
rect -1264 89 -1255 93
rect -1227 89 -1219 93
rect -1264 83 -1261 89
rect -1350 74 -1346 80
rect -1300 74 -1296 80
rect -1193 74 -1190 105
rect -1185 97 -1181 119
rect -1165 105 -1161 139
rect -1158 109 -1155 115
rect -1158 105 -1149 109
rect -1185 93 -1165 97
rect -1158 93 -1155 105
rect -1121 101 -1117 131
rect -1073 109 -1070 170
rect -1093 105 -1070 109
rect -1129 97 -1117 101
rect -1121 93 -1117 97
rect -1158 89 -1149 93
rect -1121 89 -1113 93
rect -1158 83 -1155 89
rect -1073 74 -1070 105
rect -1678 71 -1070 74
rect -1534 16 -1260 19
rect -1534 13 -1531 16
rect -1264 13 -1260 16
rect -1708 10 -1482 13
rect -1708 -163 -1705 10
rect -1591 -19 -1588 10
rect -1485 -1 -1482 10
rect -1264 10 -1155 13
rect -1448 5 -1312 9
rect -1485 -5 -1476 -1
rect -1554 -9 -1492 -5
rect -1591 -23 -1582 -19
rect -1695 -27 -1598 -23
rect -1684 -45 -1664 -41
rect -1678 -51 -1674 -45
rect -1670 -78 -1666 -71
rect -1653 -78 -1650 -36
rect -1695 -82 -1677 -78
rect -1670 -82 -1650 -78
rect -1643 -78 -1639 -27
rect -1628 -45 -1614 -41
rect -1627 -51 -1623 -45
rect -1619 -78 -1615 -71
rect -1602 -74 -1598 -31
rect -1591 -35 -1588 -23
rect -1554 -27 -1550 -9
rect -1520 -19 -1517 -13
rect -1526 -23 -1517 -19
rect -1562 -31 -1550 -27
rect -1554 -35 -1550 -31
rect -1591 -39 -1582 -35
rect -1554 -39 -1546 -35
rect -1591 -42 -1588 -39
rect -1520 -41 -1517 -23
rect -1485 -17 -1482 -5
rect -1448 -9 -1444 5
rect -1420 -5 -1418 -1
rect -1456 -13 -1444 -9
rect -1448 -17 -1444 -13
rect -1492 -24 -1489 -17
rect -1485 -21 -1476 -17
rect -1448 -21 -1440 -17
rect -1485 -27 -1482 -21
rect -1410 -32 -1406 5
rect -1492 -36 -1406 -32
rect -1554 -56 -1508 -52
rect -1591 -66 -1588 -63
rect -1591 -70 -1582 -66
rect -1643 -82 -1626 -78
rect -1619 -82 -1598 -78
rect -1591 -82 -1588 -70
rect -1554 -74 -1550 -56
rect -1520 -66 -1517 -64
rect -1526 -70 -1517 -66
rect -1562 -78 -1550 -74
rect -1554 -82 -1550 -78
rect -1670 -85 -1666 -82
rect -1619 -85 -1615 -82
rect -1591 -86 -1582 -82
rect -1554 -86 -1546 -82
rect -1591 -92 -1588 -86
rect -1678 -101 -1674 -95
rect -1627 -101 -1623 -95
rect -1520 -101 -1517 -70
rect -1512 -78 -1508 -56
rect -1492 -70 -1488 -36
rect -1485 -66 -1482 -60
rect -1485 -70 -1476 -66
rect -1512 -82 -1492 -78
rect -1485 -82 -1482 -70
rect -1448 -74 -1444 -44
rect -1400 -66 -1397 -5
rect -1316 -23 -1312 5
rect -1264 -19 -1261 10
rect -1158 -1 -1155 10
rect -1019 9 -1015 535
rect -899 517 -895 535
rect -888 531 -879 535
rect -851 531 -843 535
rect -808 521 -804 554
rect -797 565 -788 569
rect -760 565 -752 569
rect -797 556 -793 565
rect -797 552 -748 556
rect -797 529 -793 552
rect -721 547 -717 588
rect -702 556 -698 599
rect -664 555 -614 559
rect -701 547 -692 551
rect -721 543 -708 547
rect -721 536 -708 539
rect -760 535 -708 536
rect -701 535 -698 547
rect -664 543 -660 555
rect -636 547 -632 551
rect -672 539 -660 543
rect -664 535 -660 539
rect -760 532 -717 535
rect -797 525 -788 529
rect -899 513 -804 517
rect -797 513 -794 525
rect -760 521 -756 532
rect -701 531 -692 535
rect -664 531 -656 535
rect -732 525 -722 529
rect -768 517 -756 521
rect -760 513 -756 517
rect -797 509 -788 513
rect -760 509 -752 513
rect -726 506 -722 525
rect -632 506 -628 547
rect -586 506 -582 611
rect -794 502 -582 506
rect -900 228 -698 231
rect -900 214 -896 228
rect -797 222 -793 228
rect -863 217 -812 221
rect -900 210 -891 214
rect -958 206 -907 210
rect -1121 5 -1015 9
rect -1003 198 -907 202
rect -900 198 -897 210
rect -863 206 -859 217
rect -835 210 -827 214
rect -871 202 -859 206
rect -863 198 -859 202
rect -1003 92 -999 198
rect -900 194 -891 198
rect -863 194 -855 198
rect -831 176 -827 210
rect -816 195 -812 217
rect -789 195 -785 202
rect -816 191 -796 195
rect -789 191 -614 195
rect -789 188 -785 191
rect -797 176 -793 178
rect -831 172 -793 176
rect -813 168 -809 172
rect -586 168 -582 502
rect -813 164 -582 168
rect -889 152 -698 156
rect -760 141 -717 145
rect -797 134 -788 138
rect -899 130 -804 134
rect -899 100 -895 130
rect -808 111 -804 126
rect -797 122 -794 134
rect -760 130 -756 141
rect -732 134 -729 138
rect -768 126 -756 130
rect -760 122 -756 126
rect -851 107 -804 111
rect -888 100 -879 104
rect -958 96 -895 100
rect -1003 88 -895 92
rect -888 88 -885 100
rect -851 96 -847 107
rect -823 100 -819 104
rect -859 92 -847 96
rect -851 88 -847 92
rect -1158 -5 -1149 -1
rect -1227 -9 -1165 -5
rect -1264 -23 -1255 -19
rect -1316 -27 -1271 -23
rect -1356 -45 -1332 -41
rect -1420 -70 -1397 -66
rect -1456 -78 -1444 -74
rect -1448 -82 -1444 -78
rect -1485 -86 -1476 -82
rect -1448 -86 -1440 -82
rect -1485 -92 -1482 -86
rect -1400 -101 -1397 -70
rect -1350 -51 -1346 -45
rect -1342 -78 -1338 -71
rect -1326 -78 -1321 -36
rect -1361 -82 -1349 -78
rect -1342 -82 -1321 -78
rect -1316 -78 -1312 -27
rect -1301 -45 -1287 -41
rect -1300 -51 -1296 -45
rect -1292 -78 -1288 -71
rect -1275 -74 -1271 -31
rect -1264 -35 -1261 -23
rect -1227 -27 -1223 -9
rect -1193 -19 -1190 -13
rect -1199 -23 -1190 -19
rect -1235 -31 -1223 -27
rect -1227 -35 -1223 -31
rect -1264 -39 -1255 -35
rect -1227 -39 -1219 -35
rect -1264 -42 -1261 -39
rect -1193 -41 -1190 -23
rect -1158 -17 -1155 -5
rect -1121 -9 -1117 5
rect -1093 -5 -1091 -1
rect -1129 -13 -1117 -9
rect -1121 -17 -1117 -13
rect -1165 -24 -1162 -17
rect -1158 -21 -1149 -17
rect -1121 -21 -1113 -17
rect -1158 -27 -1155 -21
rect -1083 -32 -1079 5
rect -1165 -36 -1079 -32
rect -1227 -56 -1181 -52
rect -1264 -66 -1261 -63
rect -1264 -70 -1255 -66
rect -1316 -82 -1299 -78
rect -1292 -82 -1271 -78
rect -1264 -82 -1261 -70
rect -1227 -74 -1223 -56
rect -1193 -66 -1190 -64
rect -1199 -70 -1190 -66
rect -1235 -78 -1223 -74
rect -1227 -82 -1223 -78
rect -1342 -85 -1338 -82
rect -1292 -85 -1288 -82
rect -1264 -86 -1255 -82
rect -1227 -86 -1219 -82
rect -1264 -92 -1261 -86
rect -1350 -101 -1346 -95
rect -1300 -101 -1296 -95
rect -1193 -101 -1190 -70
rect -1185 -78 -1181 -56
rect -1165 -70 -1161 -36
rect -1158 -66 -1155 -60
rect -1158 -70 -1149 -66
rect -1185 -82 -1165 -78
rect -1158 -82 -1155 -70
rect -1121 -74 -1117 -44
rect -1073 -66 -1070 -5
rect -1093 -70 -1070 -66
rect -1129 -78 -1117 -74
rect -1121 -82 -1117 -78
rect -1158 -86 -1149 -82
rect -1121 -86 -1113 -82
rect -1158 -92 -1155 -86
rect -1073 -101 -1070 -70
rect -1678 -104 -1070 -101
rect -1534 -160 -1260 -157
rect -1534 -163 -1531 -160
rect -1264 -163 -1260 -160
rect -1708 -166 -1482 -163
rect -1708 -338 -1705 -166
rect -1591 -195 -1588 -166
rect -1485 -177 -1482 -166
rect -1264 -166 -1155 -163
rect -1448 -171 -1312 -167
rect -1485 -181 -1476 -177
rect -1554 -185 -1492 -181
rect -1591 -199 -1582 -195
rect -1695 -203 -1598 -199
rect -1684 -221 -1664 -217
rect -1678 -227 -1674 -221
rect -1670 -254 -1666 -247
rect -1653 -254 -1650 -212
rect -1695 -258 -1677 -254
rect -1670 -258 -1650 -254
rect -1643 -254 -1639 -203
rect -1628 -221 -1614 -217
rect -1627 -227 -1623 -221
rect -1619 -254 -1615 -247
rect -1602 -250 -1598 -207
rect -1591 -211 -1588 -199
rect -1554 -203 -1550 -185
rect -1520 -195 -1517 -189
rect -1526 -199 -1517 -195
rect -1562 -207 -1550 -203
rect -1554 -211 -1550 -207
rect -1591 -215 -1582 -211
rect -1554 -215 -1546 -211
rect -1591 -218 -1588 -215
rect -1520 -217 -1517 -199
rect -1485 -193 -1482 -181
rect -1448 -185 -1444 -171
rect -1420 -181 -1418 -177
rect -1456 -189 -1444 -185
rect -1448 -193 -1444 -189
rect -1492 -200 -1489 -193
rect -1485 -197 -1476 -193
rect -1448 -197 -1440 -193
rect -1485 -203 -1482 -197
rect -1410 -208 -1406 -171
rect -1492 -212 -1406 -208
rect -1554 -232 -1508 -228
rect -1591 -242 -1588 -239
rect -1591 -246 -1582 -242
rect -1643 -258 -1626 -254
rect -1619 -258 -1598 -254
rect -1591 -258 -1588 -246
rect -1554 -250 -1550 -232
rect -1520 -242 -1517 -240
rect -1526 -246 -1517 -242
rect -1562 -254 -1550 -250
rect -1554 -258 -1550 -254
rect -1670 -261 -1666 -258
rect -1619 -261 -1615 -258
rect -1591 -262 -1582 -258
rect -1554 -262 -1546 -258
rect -1591 -268 -1588 -262
rect -1678 -277 -1674 -271
rect -1627 -277 -1623 -271
rect -1520 -277 -1517 -246
rect -1512 -254 -1508 -232
rect -1492 -246 -1488 -212
rect -1485 -242 -1482 -236
rect -1485 -246 -1476 -242
rect -1512 -258 -1492 -254
rect -1485 -258 -1482 -246
rect -1448 -250 -1444 -220
rect -1400 -242 -1397 -181
rect -1316 -199 -1312 -171
rect -1264 -195 -1261 -166
rect -1158 -177 -1155 -166
rect -1003 -167 -999 88
rect -899 70 -895 88
rect -888 84 -879 88
rect -851 84 -843 88
rect -808 74 -804 107
rect -797 118 -788 122
rect -760 118 -752 122
rect -797 109 -793 118
rect -797 105 -748 109
rect -797 82 -793 105
rect -721 100 -717 141
rect -702 109 -698 152
rect -664 108 -614 112
rect -701 100 -692 104
rect -721 96 -708 100
rect -721 89 -708 92
rect -760 88 -708 89
rect -701 88 -698 100
rect -664 96 -660 108
rect -636 100 -632 104
rect -672 92 -660 96
rect -664 88 -660 92
rect -760 85 -717 88
rect -797 78 -788 82
rect -899 66 -804 70
rect -797 66 -794 78
rect -760 74 -756 85
rect -701 84 -692 88
rect -664 84 -656 88
rect -732 78 -722 82
rect -768 70 -756 74
rect -760 66 -756 70
rect -797 62 -788 66
rect -760 62 -752 66
rect -726 59 -722 78
rect -632 59 -628 100
rect -586 59 -582 164
rect -794 55 -582 59
rect -1121 -171 -999 -167
rect -1158 -181 -1149 -177
rect -1227 -185 -1165 -181
rect -1264 -199 -1255 -195
rect -1316 -203 -1271 -199
rect -1356 -221 -1332 -217
rect -1420 -246 -1397 -242
rect -1456 -254 -1444 -250
rect -1448 -258 -1444 -254
rect -1485 -262 -1476 -258
rect -1448 -262 -1440 -258
rect -1485 -268 -1482 -262
rect -1400 -277 -1397 -246
rect -1350 -227 -1346 -221
rect -1342 -254 -1338 -247
rect -1326 -254 -1321 -212
rect -1361 -258 -1349 -254
rect -1342 -258 -1321 -254
rect -1316 -254 -1312 -203
rect -1301 -221 -1287 -217
rect -1300 -227 -1296 -221
rect -1292 -254 -1288 -247
rect -1275 -250 -1271 -207
rect -1264 -211 -1261 -199
rect -1227 -203 -1223 -185
rect -1193 -195 -1190 -189
rect -1199 -199 -1190 -195
rect -1235 -207 -1223 -203
rect -1227 -211 -1223 -207
rect -1264 -215 -1255 -211
rect -1227 -215 -1219 -211
rect -1264 -218 -1261 -215
rect -1193 -217 -1190 -199
rect -1158 -193 -1155 -181
rect -1121 -185 -1117 -171
rect -1093 -181 -1091 -177
rect -1129 -189 -1117 -185
rect -1121 -193 -1117 -189
rect -1165 -200 -1162 -193
rect -1158 -197 -1149 -193
rect -1121 -197 -1113 -193
rect -1158 -203 -1155 -197
rect -1083 -208 -1079 -171
rect -1165 -212 -1079 -208
rect -1227 -232 -1181 -228
rect -1264 -242 -1261 -239
rect -1264 -246 -1255 -242
rect -1316 -258 -1299 -254
rect -1292 -258 -1271 -254
rect -1264 -258 -1261 -246
rect -1227 -250 -1223 -232
rect -1193 -242 -1190 -240
rect -1199 -246 -1190 -242
rect -1235 -254 -1223 -250
rect -1227 -258 -1223 -254
rect -1342 -261 -1338 -258
rect -1292 -261 -1288 -258
rect -1264 -262 -1255 -258
rect -1227 -262 -1219 -258
rect -1264 -268 -1261 -262
rect -1350 -277 -1346 -271
rect -1300 -277 -1296 -271
rect -1193 -277 -1190 -246
rect -1185 -254 -1181 -232
rect -1165 -246 -1161 -212
rect -1158 -242 -1155 -236
rect -1158 -246 -1149 -242
rect -1185 -258 -1165 -254
rect -1158 -258 -1155 -246
rect -1121 -250 -1117 -220
rect -1073 -242 -1070 -181
rect -1093 -246 -1070 -242
rect -1129 -254 -1117 -250
rect -1121 -258 -1117 -254
rect -1158 -262 -1149 -258
rect -1121 -262 -1113 -258
rect -1158 -268 -1155 -262
rect -1073 -277 -1070 -246
rect -1678 -280 -1070 -277
rect -900 -275 -698 -272
rect -900 -289 -896 -275
rect -797 -281 -793 -275
rect -863 -286 -812 -282
rect -900 -293 -891 -289
rect -969 -297 -907 -293
rect -998 -305 -907 -301
rect -900 -305 -897 -293
rect -863 -297 -859 -286
rect -835 -293 -827 -289
rect -871 -301 -859 -297
rect -863 -305 -859 -301
rect -1534 -335 -1260 -332
rect -1534 -338 -1531 -335
rect -1264 -338 -1260 -335
rect -1708 -341 -1482 -338
rect -1591 -370 -1588 -341
rect -1485 -352 -1482 -341
rect -1264 -341 -1155 -338
rect -1448 -346 -1312 -342
rect -1485 -356 -1476 -352
rect -1554 -360 -1492 -356
rect -1591 -374 -1582 -370
rect -1712 -378 -1598 -374
rect -1684 -396 -1664 -392
rect -1678 -402 -1674 -396
rect -1670 -429 -1666 -422
rect -1653 -429 -1650 -387
rect -1712 -433 -1677 -429
rect -1670 -433 -1650 -429
rect -1643 -429 -1639 -378
rect -1628 -396 -1614 -392
rect -1627 -402 -1623 -396
rect -1619 -429 -1615 -422
rect -1602 -425 -1598 -382
rect -1591 -386 -1588 -374
rect -1554 -378 -1550 -360
rect -1520 -370 -1517 -364
rect -1526 -374 -1517 -370
rect -1562 -382 -1550 -378
rect -1554 -386 -1550 -382
rect -1591 -390 -1582 -386
rect -1554 -390 -1546 -386
rect -1591 -393 -1588 -390
rect -1520 -392 -1517 -374
rect -1485 -368 -1482 -356
rect -1448 -360 -1444 -346
rect -1420 -356 -1418 -352
rect -1456 -364 -1444 -360
rect -1448 -368 -1444 -364
rect -1492 -375 -1489 -368
rect -1485 -372 -1476 -368
rect -1448 -372 -1440 -368
rect -1485 -378 -1482 -372
rect -1410 -383 -1406 -346
rect -1492 -387 -1406 -383
rect -1554 -407 -1508 -403
rect -1591 -417 -1588 -414
rect -1591 -421 -1582 -417
rect -1643 -433 -1626 -429
rect -1619 -433 -1598 -429
rect -1591 -433 -1588 -421
rect -1554 -425 -1550 -407
rect -1520 -417 -1517 -415
rect -1526 -421 -1517 -417
rect -1562 -429 -1550 -425
rect -1554 -433 -1550 -429
rect -1670 -436 -1666 -433
rect -1619 -436 -1615 -433
rect -1591 -437 -1582 -433
rect -1554 -437 -1546 -433
rect -1591 -443 -1588 -437
rect -1678 -452 -1674 -446
rect -1627 -452 -1623 -446
rect -1520 -452 -1517 -421
rect -1512 -429 -1508 -407
rect -1492 -421 -1488 -387
rect -1485 -417 -1482 -411
rect -1485 -421 -1476 -417
rect -1512 -433 -1492 -429
rect -1485 -433 -1482 -421
rect -1448 -425 -1444 -395
rect -1400 -417 -1397 -356
rect -1316 -374 -1312 -346
rect -1264 -370 -1261 -341
rect -1158 -352 -1155 -341
rect -998 -342 -994 -305
rect -900 -309 -891 -305
rect -863 -309 -855 -305
rect -831 -327 -827 -293
rect -816 -308 -812 -286
rect -789 -308 -785 -301
rect -816 -312 -796 -308
rect -789 -312 -614 -308
rect -789 -315 -785 -312
rect -797 -327 -793 -325
rect -831 -331 -793 -327
rect -815 -335 -811 -331
rect -586 -335 -582 55
rect -815 -339 -582 -335
rect -1121 -346 -994 -342
rect -1158 -356 -1149 -352
rect -1227 -360 -1165 -356
rect -1264 -374 -1255 -370
rect -1316 -378 -1271 -374
rect -1356 -396 -1332 -392
rect -1420 -421 -1397 -417
rect -1456 -429 -1444 -425
rect -1448 -433 -1444 -429
rect -1485 -437 -1476 -433
rect -1448 -437 -1440 -433
rect -1485 -443 -1482 -437
rect -1400 -452 -1397 -421
rect -1350 -402 -1346 -396
rect -1342 -429 -1338 -422
rect -1326 -429 -1321 -387
rect -1361 -433 -1349 -429
rect -1342 -433 -1321 -429
rect -1316 -429 -1312 -378
rect -1301 -396 -1287 -392
rect -1300 -402 -1296 -396
rect -1292 -429 -1288 -422
rect -1275 -425 -1271 -382
rect -1264 -386 -1261 -374
rect -1227 -378 -1223 -360
rect -1193 -370 -1190 -364
rect -1199 -374 -1190 -370
rect -1235 -382 -1223 -378
rect -1227 -386 -1223 -382
rect -1264 -390 -1255 -386
rect -1227 -390 -1219 -386
rect -1264 -393 -1261 -390
rect -1193 -392 -1190 -374
rect -1158 -368 -1155 -356
rect -1121 -360 -1117 -346
rect -1093 -356 -1091 -352
rect -1129 -364 -1117 -360
rect -1121 -368 -1117 -364
rect -1165 -375 -1162 -368
rect -1158 -372 -1149 -368
rect -1121 -372 -1113 -368
rect -1158 -378 -1155 -372
rect -1083 -383 -1079 -346
rect -1165 -387 -1079 -383
rect -1227 -407 -1181 -403
rect -1264 -417 -1261 -414
rect -1264 -421 -1255 -417
rect -1316 -433 -1299 -429
rect -1292 -433 -1271 -429
rect -1264 -433 -1261 -421
rect -1227 -425 -1223 -407
rect -1193 -417 -1190 -415
rect -1199 -421 -1190 -417
rect -1235 -429 -1223 -425
rect -1227 -433 -1223 -429
rect -1342 -436 -1338 -433
rect -1292 -436 -1288 -433
rect -1264 -437 -1255 -433
rect -1227 -437 -1219 -433
rect -1264 -443 -1261 -437
rect -1350 -452 -1346 -446
rect -1300 -452 -1296 -446
rect -1193 -452 -1190 -421
rect -1185 -429 -1181 -407
rect -1165 -421 -1161 -387
rect -1158 -417 -1155 -411
rect -1158 -421 -1149 -417
rect -1185 -433 -1165 -429
rect -1158 -433 -1155 -421
rect -1121 -425 -1117 -395
rect -1073 -417 -1070 -356
rect -998 -411 -994 -346
rect -889 -351 -698 -347
rect -760 -362 -717 -358
rect -797 -369 -788 -365
rect -899 -373 -804 -369
rect -899 -403 -895 -373
rect -808 -392 -804 -377
rect -797 -381 -794 -369
rect -760 -373 -756 -362
rect -732 -369 -729 -365
rect -768 -377 -756 -373
rect -760 -381 -756 -377
rect -851 -396 -804 -392
rect -888 -403 -879 -399
rect -969 -407 -895 -403
rect -998 -415 -895 -411
rect -888 -415 -885 -403
rect -851 -407 -847 -396
rect -823 -403 -819 -399
rect -859 -411 -847 -407
rect -851 -415 -847 -411
rect -1093 -421 -1070 -417
rect -1129 -429 -1117 -425
rect -1121 -433 -1117 -429
rect -1158 -437 -1149 -433
rect -1121 -437 -1113 -433
rect -1158 -443 -1155 -437
rect -1073 -452 -1070 -421
rect -899 -433 -895 -415
rect -888 -419 -879 -415
rect -851 -419 -843 -415
rect -808 -429 -804 -396
rect -797 -385 -788 -381
rect -760 -385 -752 -381
rect -797 -394 -793 -385
rect -797 -398 -748 -394
rect -797 -421 -793 -398
rect -721 -403 -717 -362
rect -702 -394 -698 -351
rect -664 -395 -614 -391
rect -701 -403 -692 -399
rect -721 -407 -708 -403
rect -721 -414 -708 -411
rect -760 -415 -708 -414
rect -701 -415 -698 -403
rect -664 -407 -660 -395
rect -636 -403 -632 -399
rect -672 -411 -660 -407
rect -664 -415 -660 -411
rect -760 -418 -717 -415
rect -797 -425 -788 -421
rect -899 -437 -804 -433
rect -797 -437 -794 -425
rect -760 -429 -756 -418
rect -701 -419 -692 -415
rect -664 -419 -656 -415
rect -732 -425 -722 -421
rect -768 -433 -756 -429
rect -760 -437 -756 -433
rect -797 -441 -788 -437
rect -760 -441 -752 -437
rect -726 -444 -722 -425
rect -632 -444 -628 -403
rect -586 -444 -582 -339
rect -794 -448 -582 -444
rect -1723 -455 -1070 -452
rect -1723 -462 -1720 -455
rect -585 -462 -582 -448
rect -1723 -465 -582 -462
rect -1723 -518 -1720 -465
rect -567 -500 -563 862
rect -454 852 -451 862
rect -356 859 -352 862
rect -422 855 -362 858
rect -422 852 -419 855
rect -477 848 -473 852
rect -454 848 -448 852
rect -423 848 -416 852
rect -540 832 -536 847
rect -477 844 -461 848
rect -465 836 -461 840
rect -454 836 -451 848
rect -423 844 -419 848
rect -428 840 -419 844
rect -454 832 -448 836
rect -540 828 -461 832
rect -540 769 -536 828
rect -502 791 -498 819
rect -487 820 -461 824
rect -454 820 -451 832
rect -423 828 -419 840
rect -428 824 -419 828
rect -373 820 -370 852
rect -365 830 -362 855
rect -348 830 -344 839
rect -365 826 -355 830
rect -348 826 -338 830
rect -348 823 -344 826
rect -540 765 -502 769
rect -487 759 -483 820
rect -454 816 -448 820
rect -376 816 -370 820
rect -454 813 -451 816
rect -373 810 -370 816
rect -356 810 -352 813
rect -462 807 -344 810
rect -323 795 -320 862
rect -452 792 -320 795
rect -469 772 -459 775
rect -452 771 -449 792
rect -364 789 -360 792
rect -420 782 -370 785
rect -420 779 -417 782
rect -426 775 -414 779
rect -452 767 -446 771
rect -473 763 -459 767
rect -487 755 -459 759
rect -452 755 -449 767
rect -421 763 -417 775
rect -426 759 -417 763
rect -381 755 -378 779
rect -373 760 -370 782
rect -356 760 -352 769
rect -373 756 -363 760
rect -356 756 -333 760
rect -487 681 -483 755
rect -452 751 -446 755
rect -384 751 -378 755
rect -356 753 -352 756
rect -381 740 -378 751
rect -364 740 -360 743
rect -381 737 -352 740
rect -323 720 -320 792
rect -452 717 -320 720
rect -452 693 -449 717
rect -373 714 -369 717
rect -420 696 -380 700
rect -420 693 -416 696
rect -452 689 -446 693
rect -420 689 -413 693
rect -470 685 -459 689
rect -487 677 -459 681
rect -452 677 -449 689
rect -420 685 -416 689
rect -384 685 -380 696
rect -365 685 -361 694
rect -426 681 -416 685
rect -384 681 -372 685
rect -365 681 -319 685
rect -365 678 -361 681
rect -548 630 -528 651
rect -487 607 -483 677
rect -452 673 -446 677
rect -393 673 -387 677
rect -390 665 -387 673
rect -373 665 -369 668
rect -390 662 -369 665
rect -305 644 -302 947
rect -64 919 -60 1066
rect -93 898 169 902
rect -93 863 -89 898
rect -244 860 -86 863
rect -280 843 -240 847
rect -280 830 -276 843
rect -267 835 -240 839
rect -267 761 -263 835
rect -288 757 -263 761
rect -256 827 -240 831
rect -256 685 -252 827
rect -280 681 -252 685
rect -246 819 -240 823
rect -233 819 -230 860
rect -142 854 -110 857
rect -142 851 -139 854
rect -147 847 -139 851
rect -125 847 -119 851
rect -143 843 -139 847
rect -143 839 -135 843
rect -143 827 -139 839
rect -122 835 -119 847
rect -125 831 -119 835
rect -143 823 -135 827
rect -122 819 -119 831
rect -113 827 -110 854
rect -104 856 -100 860
rect -65 846 -61 889
rect 107 887 150 891
rect 70 880 79 884
rect -32 876 63 880
rect -32 846 -28 876
rect 59 857 63 872
rect 70 868 73 880
rect 107 876 111 887
rect 135 880 138 884
rect 99 872 111 876
rect 107 868 111 872
rect 16 853 63 857
rect -21 846 -12 850
rect -65 842 -28 846
rect -96 827 -92 836
rect -54 834 -28 838
rect -21 834 -18 846
rect 16 842 20 853
rect 44 846 48 850
rect 8 838 20 842
rect 16 834 20 838
rect -113 823 -103 827
rect -96 823 -86 827
rect -96 820 -92 823
rect -470 641 -302 644
rect -246 629 -243 819
rect -233 815 -227 819
rect -125 815 -119 819
rect -122 807 -119 815
rect -54 820 -50 834
rect -32 816 -28 834
rect -21 830 -12 834
rect 16 830 24 834
rect 59 820 63 853
rect 70 864 79 868
rect 107 864 115 868
rect 70 855 74 864
rect 70 851 119 855
rect 70 828 74 851
rect 146 846 150 887
rect 165 855 169 898
rect 249 858 269 867
rect 203 854 269 858
rect 166 846 175 850
rect 146 842 159 846
rect 146 835 159 838
rect 107 834 159 835
rect 166 834 169 846
rect 203 842 207 854
rect 231 846 235 850
rect 249 846 269 854
rect 195 838 207 842
rect 203 834 207 838
rect 107 831 150 834
rect 70 824 79 828
rect -32 812 63 816
rect 70 812 73 824
rect 107 820 111 831
rect 166 830 175 834
rect 203 830 211 834
rect 135 824 145 828
rect 99 816 111 820
rect 107 812 111 816
rect -104 807 -100 810
rect 70 808 79 812
rect 107 808 115 812
rect -122 805 -40 807
rect 141 805 145 824
rect 235 805 239 846
rect -122 804 239 805
rect -44 801 239 804
rect -54 774 -50 794
rect -475 626 -243 629
rect -229 770 -50 774
rect -229 607 -225 770
rect -487 603 -225 607
rect -548 559 -528 568
rect -487 559 -483 603
rect -548 555 -483 559
rect -548 547 -528 555
rect -548 184 -528 205
rect -548 101 -528 122
rect -548 -319 -528 -298
rect -548 -402 -528 -381
rect -1708 -503 -563 -500
rect -1708 -518 -1705 -503
<< m2contact >>
rect -1708 1543 -1703 1548
rect -1501 1540 -1496 1545
rect -1653 1499 -1648 1504
rect -1663 1490 -1658 1495
rect -1606 1499 -1601 1504
rect -1632 1490 -1627 1495
rect -1613 1490 -1608 1495
rect -1417 1530 -1412 1535
rect -1493 1506 -1488 1511
rect -1448 1506 -1442 1511
rect -1400 1530 -1395 1535
rect -1592 1488 -1587 1493
rect -1520 1489 -1515 1494
rect -1592 1472 -1587 1477
rect -1519 1471 -1514 1476
rect -1751 1330 -1746 1335
rect -1751 1155 -1746 1160
rect -1751 980 -1746 985
rect -1751 804 -1746 809
rect -1751 629 -1746 634
rect -1751 323 -1746 328
rect -1751 148 -1746 153
rect -1751 -27 -1746 -22
rect -1751 -203 -1746 -198
rect -1751 -378 -1746 -373
rect -1448 1491 -1442 1496
rect -1484 1475 -1479 1480
rect -1268 1522 -1263 1528
rect -1174 1540 -1169 1545
rect -1325 1499 -1320 1504
rect -1343 1494 -1338 1499
rect -1365 1452 -1360 1457
rect -1279 1499 -1274 1504
rect -1305 1490 -1300 1495
rect -1286 1490 -1281 1495
rect -1090 1530 -1085 1535
rect -1166 1506 -1161 1511
rect -1121 1506 -1115 1511
rect -1073 1530 -1068 1535
rect -1265 1488 -1260 1493
rect -1193 1489 -1188 1494
rect -1265 1472 -1260 1477
rect -1192 1471 -1187 1476
rect -1121 1491 -1115 1496
rect -1157 1475 -1152 1480
rect -1734 1275 -1729 1280
rect -1734 1100 -1729 1105
rect -1734 925 -1729 930
rect -1734 749 -1729 754
rect -1734 573 -1729 578
rect -1709 1412 -1704 1417
rect -694 1398 -689 1403
rect -1720 1252 -1715 1257
rect -1501 1362 -1496 1367
rect -1699 1330 -1694 1335
rect -1653 1321 -1648 1326
rect -1663 1312 -1658 1317
rect -1699 1275 -1694 1280
rect -1606 1321 -1601 1326
rect -1632 1312 -1627 1317
rect -1613 1312 -1608 1317
rect -1417 1352 -1412 1357
rect -1493 1328 -1488 1333
rect -1448 1328 -1442 1333
rect -1400 1352 -1395 1357
rect -1592 1310 -1587 1315
rect -1520 1311 -1515 1316
rect -1592 1294 -1587 1299
rect -1519 1293 -1514 1298
rect -1682 1252 -1677 1257
rect -1448 1313 -1442 1318
rect -1484 1297 -1479 1302
rect -1268 1344 -1263 1350
rect -1174 1362 -1169 1367
rect -1325 1321 -1320 1326
rect -1343 1316 -1338 1321
rect -1365 1274 -1360 1279
rect -1279 1321 -1274 1326
rect -1305 1312 -1300 1317
rect -1286 1312 -1281 1317
rect -1090 1352 -1085 1357
rect -1166 1328 -1161 1333
rect -1121 1328 -1115 1333
rect -1073 1352 -1068 1357
rect -1265 1310 -1260 1315
rect -1193 1311 -1188 1316
rect -1265 1294 -1260 1299
rect -1192 1293 -1187 1298
rect -1121 1313 -1115 1318
rect -1157 1297 -1152 1302
rect -1056 1273 -1051 1278
rect -614 1362 -609 1367
rect -582 1450 -577 1455
rect -572 1398 -567 1403
rect -885 1318 -880 1323
rect -917 1273 -912 1278
rect -725 1304 -720 1309
rect -885 1275 -880 1280
rect -815 1270 -810 1275
rect -1720 1077 -1715 1082
rect -1502 1187 -1497 1192
rect -1700 1155 -1695 1160
rect -1654 1146 -1649 1151
rect -1664 1137 -1659 1142
rect -1700 1100 -1695 1105
rect -1607 1146 -1602 1151
rect -1633 1137 -1628 1142
rect -1614 1137 -1609 1142
rect -1418 1177 -1413 1182
rect -1494 1153 -1489 1158
rect -1449 1153 -1443 1158
rect -1401 1177 -1396 1182
rect -1593 1135 -1588 1140
rect -1521 1136 -1516 1141
rect -1593 1119 -1588 1124
rect -1520 1118 -1515 1123
rect -1683 1077 -1678 1082
rect -1449 1138 -1443 1143
rect -1485 1122 -1480 1127
rect -1269 1169 -1264 1175
rect -1175 1187 -1170 1192
rect -1326 1146 -1321 1151
rect -1344 1141 -1339 1146
rect -1366 1099 -1361 1104
rect -1280 1146 -1275 1151
rect -1306 1137 -1301 1142
rect -1287 1137 -1282 1142
rect -1091 1177 -1086 1182
rect -1167 1153 -1162 1158
rect -1122 1153 -1116 1158
rect -1061 1186 -1056 1191
rect -1074 1177 -1069 1182
rect -1266 1135 -1261 1140
rect -1194 1136 -1189 1141
rect -1266 1119 -1261 1124
rect -1193 1118 -1188 1123
rect -1122 1138 -1116 1143
rect -1158 1122 -1153 1127
rect -1720 902 -1715 907
rect -1502 1012 -1497 1017
rect -1700 980 -1695 985
rect -1654 971 -1649 976
rect -1664 962 -1659 967
rect -1700 925 -1695 930
rect -1607 971 -1602 976
rect -1633 962 -1628 967
rect -1614 962 -1609 967
rect -1418 1002 -1413 1007
rect -1494 978 -1489 983
rect -1449 978 -1443 983
rect -1401 1002 -1396 1007
rect -1593 960 -1588 965
rect -1521 961 -1516 966
rect -1593 944 -1588 949
rect -1520 943 -1515 948
rect -1683 902 -1678 907
rect -1449 963 -1443 968
rect -1485 947 -1480 952
rect -1269 994 -1264 1000
rect -1175 1012 -1170 1017
rect -1063 1012 -1058 1017
rect -1326 971 -1321 976
rect -1344 966 -1339 971
rect -1366 924 -1361 929
rect -1280 971 -1275 976
rect -1306 962 -1301 967
rect -1287 962 -1282 967
rect -1091 1002 -1086 1007
rect -1167 978 -1162 983
rect -1122 978 -1116 983
rect -1074 1002 -1069 1007
rect -1266 960 -1261 965
rect -1194 961 -1189 966
rect -1266 944 -1261 949
rect -1193 943 -1188 948
rect -1122 963 -1116 968
rect -1158 947 -1153 952
rect -1720 726 -1715 731
rect -1502 836 -1497 841
rect -1700 804 -1695 809
rect -1654 795 -1649 800
rect -1664 786 -1659 791
rect -1700 749 -1695 754
rect -1607 795 -1602 800
rect -1633 786 -1628 791
rect -1614 786 -1609 791
rect -1418 826 -1413 831
rect -1494 802 -1489 807
rect -1449 802 -1443 807
rect -1401 826 -1396 831
rect -1593 784 -1588 789
rect -1521 785 -1516 790
rect -1593 768 -1588 773
rect -1520 767 -1515 772
rect -1683 726 -1678 731
rect -1449 787 -1443 792
rect -1485 771 -1480 776
rect -1269 818 -1264 824
rect -1175 836 -1170 841
rect -1326 795 -1321 800
rect -1344 790 -1339 795
rect -1366 748 -1361 753
rect -1280 795 -1275 800
rect -1306 786 -1301 791
rect -1287 786 -1282 791
rect -1091 826 -1086 831
rect -1167 802 -1162 807
rect -1122 802 -1116 807
rect -1062 835 -1057 840
rect -1074 826 -1069 831
rect -1266 784 -1261 789
rect -1194 785 -1189 790
rect -1266 768 -1261 773
rect -1193 767 -1188 772
rect -1122 787 -1116 792
rect -1158 771 -1153 776
rect -1710 661 -1705 666
rect -1502 661 -1497 666
rect -1717 629 -1712 634
rect -1654 620 -1649 625
rect -1664 611 -1659 616
rect -1717 573 -1712 578
rect -1607 620 -1602 625
rect -1633 611 -1628 616
rect -1614 611 -1609 616
rect -1418 651 -1413 656
rect -1494 627 -1489 632
rect -1449 627 -1443 632
rect -1401 651 -1396 656
rect -1593 609 -1588 614
rect -1521 610 -1516 615
rect -1593 593 -1588 598
rect -1520 592 -1515 597
rect -1449 612 -1443 617
rect -1485 596 -1480 601
rect -1269 643 -1264 649
rect -1175 661 -1170 666
rect -1326 620 -1321 625
rect -1344 615 -1339 620
rect -1366 573 -1361 578
rect -1280 620 -1275 625
rect -1306 611 -1301 616
rect -1287 611 -1282 616
rect -1091 651 -1086 656
rect -1167 627 -1162 632
rect -1122 627 -1116 632
rect -1067 660 -1062 665
rect -1074 651 -1069 656
rect -1266 609 -1261 614
rect -1194 610 -1189 615
rect -1266 593 -1261 598
rect -1193 592 -1188 597
rect -1122 612 -1116 617
rect -1158 596 -1153 601
rect -1734 268 -1729 273
rect -1734 93 -1729 98
rect -1734 -82 -1729 -77
rect -1734 -258 -1729 -253
rect -1734 -434 -1729 -429
rect -1709 507 -1704 512
rect -1720 245 -1715 250
rect -1501 355 -1496 360
rect -1699 323 -1694 328
rect -1653 314 -1648 319
rect -1663 305 -1658 310
rect -1699 268 -1694 273
rect -1606 314 -1601 319
rect -1632 305 -1627 310
rect -1613 305 -1608 310
rect -1417 345 -1412 350
rect -1493 321 -1488 326
rect -1448 321 -1442 326
rect -1400 345 -1395 350
rect -1592 303 -1587 308
rect -1520 304 -1515 309
rect -1592 287 -1587 292
rect -1519 286 -1514 291
rect -1682 245 -1677 250
rect -1448 306 -1442 311
rect -1484 290 -1479 295
rect -1268 337 -1263 343
rect -1174 355 -1169 360
rect -744 1276 -739 1281
rect -694 1322 -689 1327
rect -699 1275 -694 1280
rect -614 1279 -609 1284
rect -628 1271 -623 1276
rect -572 1322 -567 1327
rect -916 1186 -911 1191
rect -698 1032 -693 1037
rect -614 996 -609 1001
rect -582 1215 -577 1220
rect -582 1160 -577 1165
rect -572 1032 -567 1037
rect -889 952 -884 957
rect -933 904 -928 909
rect -729 938 -724 943
rect -889 909 -884 914
rect -819 904 -814 909
rect -1325 314 -1320 319
rect -1343 309 -1338 314
rect -1365 267 -1360 272
rect -1279 314 -1274 319
rect -1305 305 -1300 310
rect -1286 305 -1281 310
rect -1090 345 -1085 350
rect -1166 321 -1161 326
rect -1121 321 -1115 326
rect -1073 345 -1068 350
rect -1265 303 -1260 308
rect -1193 304 -1188 309
rect -1265 287 -1260 292
rect -1192 286 -1187 291
rect -1121 306 -1115 311
rect -1157 290 -1152 295
rect -1720 70 -1715 75
rect -1502 180 -1497 185
rect -1700 148 -1695 153
rect -1654 139 -1649 144
rect -1664 130 -1659 135
rect -1700 93 -1695 98
rect -1607 139 -1602 144
rect -1633 130 -1628 135
rect -1614 130 -1609 135
rect -1418 170 -1413 175
rect -1494 146 -1489 151
rect -1449 146 -1443 151
rect -1401 170 -1396 175
rect -1593 128 -1588 133
rect -1521 129 -1516 134
rect -1593 112 -1588 117
rect -1520 111 -1515 116
rect -1683 70 -1678 75
rect -1449 131 -1443 136
rect -1485 115 -1480 120
rect -1269 162 -1264 168
rect -1175 180 -1170 185
rect -748 910 -743 915
rect -698 956 -693 961
rect -703 909 -698 914
rect -614 913 -609 918
rect -632 905 -627 910
rect -572 956 -567 961
rect -698 674 -693 679
rect -949 652 -944 657
rect -614 638 -609 643
rect -525 1510 -520 1515
rect -499 1510 -494 1515
rect -553 1362 -548 1367
rect -528 1362 -523 1367
rect -499 1455 -494 1460
rect -241 1440 -236 1445
rect -381 1420 -376 1425
rect -502 1362 -497 1367
rect -361 1420 -356 1425
rect -227 1383 -222 1388
rect -221 1338 -216 1343
rect -201 1383 -196 1388
rect -158 1379 -153 1384
rect 2 1365 7 1370
rect -158 1336 -153 1341
rect -88 1331 -83 1336
rect -325 1287 -320 1292
rect -206 1288 -201 1293
rect -17 1337 -12 1342
rect 28 1336 33 1341
rect 99 1332 104 1337
rect -180 1288 -175 1293
rect -553 1279 -548 1284
rect -192 1275 -187 1280
rect -266 1268 -261 1273
rect -325 1243 -320 1248
rect -507 1215 -502 1220
rect -334 1214 -329 1219
rect -505 1160 -500 1165
rect -394 1158 -389 1163
rect -342 1158 -337 1163
rect -314 1214 -309 1219
rect -493 1147 -488 1152
rect -130 1212 -125 1217
rect -241 1167 -236 1172
rect -93 1190 -88 1195
rect 30 1198 35 1203
rect -130 1169 -125 1174
rect -342 1133 -337 1138
rect -553 996 -548 1001
rect -528 996 -523 1001
rect -553 913 -548 918
rect -416 1081 -411 1086
rect -60 1164 -55 1169
rect -121 1135 -116 1140
rect 11 1170 16 1175
rect 56 1169 61 1174
rect 127 1165 132 1170
rect -153 1119 -148 1124
rect -357 1050 -352 1055
rect -180 1026 -175 1031
rect -467 996 -462 1001
rect -159 985 -154 990
rect -117 985 -112 990
rect -540 900 -535 905
rect -582 805 -577 810
rect -572 674 -567 679
rect -889 594 -884 599
rect -729 580 -724 585
rect -889 551 -884 556
rect -949 542 -944 547
rect -819 546 -814 551
rect -1326 139 -1321 144
rect -1344 134 -1339 139
rect -1366 92 -1361 97
rect -1280 139 -1275 144
rect -1306 130 -1301 135
rect -1287 130 -1282 135
rect -1091 170 -1086 175
rect -1167 146 -1162 151
rect -1122 146 -1116 151
rect -1074 170 -1069 175
rect -1266 128 -1261 133
rect -1194 129 -1189 134
rect -1266 112 -1261 117
rect -1193 111 -1188 116
rect -1122 131 -1116 136
rect -1158 115 -1153 120
rect -1720 -105 -1715 -100
rect -1502 5 -1497 10
rect -1700 -27 -1695 -22
rect -1654 -36 -1649 -31
rect -1664 -45 -1659 -40
rect -1700 -82 -1695 -77
rect -1607 -36 -1602 -31
rect -1633 -45 -1628 -40
rect -1614 -45 -1609 -40
rect -1418 -5 -1413 0
rect -1494 -29 -1489 -24
rect -1449 -29 -1443 -24
rect -1401 -5 -1396 0
rect -1593 -47 -1588 -42
rect -1521 -46 -1516 -41
rect -1593 -63 -1588 -58
rect -1520 -64 -1515 -59
rect -1683 -105 -1678 -100
rect -1449 -44 -1443 -39
rect -1485 -60 -1480 -55
rect -1269 -13 -1264 -7
rect -1175 5 -1170 10
rect -748 552 -743 557
rect -698 598 -693 603
rect -703 551 -698 556
rect -614 555 -609 560
rect -632 547 -627 552
rect -572 598 -567 603
rect -698 227 -693 232
rect -963 205 -958 210
rect -614 191 -609 196
rect -572 227 -567 232
rect -889 147 -884 152
rect -729 133 -724 138
rect -889 104 -884 109
rect -963 95 -958 100
rect -819 99 -814 104
rect -1326 -36 -1321 -31
rect -1344 -41 -1339 -36
rect -1366 -83 -1361 -78
rect -1280 -36 -1275 -31
rect -1306 -45 -1301 -40
rect -1287 -45 -1282 -40
rect -1091 -5 -1086 0
rect -1167 -29 -1162 -24
rect -1122 -29 -1116 -24
rect -1074 -5 -1069 0
rect -1266 -47 -1261 -42
rect -1194 -46 -1189 -41
rect -1266 -63 -1261 -58
rect -1193 -64 -1188 -59
rect -1122 -44 -1116 -39
rect -1158 -60 -1153 -55
rect -1720 -281 -1715 -276
rect -1502 -171 -1497 -166
rect -1700 -203 -1695 -198
rect -1654 -212 -1649 -207
rect -1664 -221 -1659 -216
rect -1700 -258 -1695 -253
rect -1607 -212 -1602 -207
rect -1633 -221 -1628 -216
rect -1614 -221 -1609 -216
rect -1418 -181 -1413 -176
rect -1494 -205 -1489 -200
rect -1449 -205 -1443 -200
rect -1401 -181 -1396 -176
rect -1593 -223 -1588 -218
rect -1521 -222 -1516 -217
rect -1593 -239 -1588 -234
rect -1520 -240 -1515 -235
rect -1683 -281 -1678 -276
rect -1449 -220 -1443 -215
rect -1485 -236 -1480 -231
rect -1269 -189 -1264 -183
rect -1175 -171 -1170 -166
rect -748 105 -743 110
rect -698 151 -693 156
rect -703 104 -698 109
rect -614 108 -609 113
rect -632 100 -627 105
rect -572 151 -567 156
rect -1326 -212 -1321 -207
rect -1344 -217 -1339 -212
rect -1366 -259 -1361 -254
rect -1280 -212 -1275 -207
rect -1306 -221 -1301 -216
rect -1287 -221 -1282 -216
rect -1091 -181 -1086 -176
rect -1167 -205 -1162 -200
rect -1122 -205 -1116 -200
rect -1074 -181 -1069 -176
rect -1266 -223 -1261 -218
rect -1194 -222 -1189 -217
rect -1266 -239 -1261 -234
rect -1193 -240 -1188 -235
rect -1122 -220 -1116 -215
rect -1158 -236 -1153 -231
rect -698 -276 -693 -271
rect -974 -297 -969 -292
rect -1710 -346 -1705 -341
rect -1502 -346 -1497 -341
rect -1717 -378 -1712 -373
rect -1654 -387 -1649 -382
rect -1664 -396 -1659 -391
rect -1717 -434 -1712 -429
rect -1607 -387 -1602 -382
rect -1633 -396 -1628 -391
rect -1614 -396 -1609 -391
rect -1418 -356 -1413 -351
rect -1494 -380 -1489 -375
rect -1449 -380 -1443 -375
rect -1401 -356 -1396 -351
rect -1593 -398 -1588 -393
rect -1521 -397 -1516 -392
rect -1593 -414 -1588 -409
rect -1520 -415 -1515 -410
rect -1449 -395 -1443 -390
rect -1485 -411 -1480 -406
rect -1269 -364 -1264 -358
rect -1175 -346 -1170 -341
rect -614 -312 -609 -307
rect -572 -276 -567 -271
rect -1326 -387 -1321 -382
rect -1344 -392 -1339 -387
rect -1366 -434 -1361 -429
rect -1280 -387 -1275 -382
rect -1306 -396 -1301 -391
rect -1287 -396 -1282 -391
rect -1091 -356 -1086 -351
rect -1167 -380 -1162 -375
rect -1122 -380 -1116 -375
rect -1074 -356 -1069 -351
rect -1266 -398 -1261 -393
rect -1194 -397 -1189 -392
rect -1266 -414 -1261 -409
rect -1193 -415 -1188 -410
rect -1122 -395 -1116 -390
rect -1158 -411 -1153 -406
rect -889 -356 -884 -351
rect -974 -407 -969 -402
rect -729 -370 -724 -365
rect -889 -399 -884 -394
rect -819 -404 -814 -399
rect -748 -398 -743 -393
rect -698 -352 -693 -347
rect -703 -399 -698 -394
rect -614 -395 -609 -390
rect -632 -403 -627 -398
rect -572 -352 -567 -347
rect -1709 -500 -1704 -495
rect -477 852 -472 857
rect -540 847 -535 852
rect -470 836 -465 841
rect -503 819 -498 824
rect -503 786 -498 791
rect -338 825 -333 830
rect -502 764 -497 769
rect -467 805 -462 810
rect -344 805 -339 810
rect -320 860 -315 865
rect -475 772 -469 778
rect -479 762 -473 768
rect -333 756 -328 761
rect -352 735 -347 740
rect -475 684 -470 689
rect -319 680 -314 685
rect -553 638 -548 643
rect -540 625 -535 630
rect -374 657 -369 662
rect -475 640 -470 645
rect -65 914 -60 919
rect -249 859 -244 864
rect -65 889 -60 894
rect -22 893 -17 898
rect -280 825 -275 830
rect -293 756 -288 761
rect -285 680 -280 685
rect 138 879 143 884
rect -22 850 -17 855
rect 48 845 53 850
rect -480 625 -475 630
rect -127 803 -122 808
rect -54 815 -49 820
rect 119 851 124 856
rect 164 850 169 855
rect 235 846 240 851
rect -54 794 -49 799
rect -553 555 -548 560
rect -553 191 -548 196
rect -553 108 -548 113
rect -553 -312 -548 -307
rect -553 -395 -548 -390
<< metal2 >>
rect -1618 1555 -1361 1558
rect -1708 1417 -1705 1543
rect -1618 1503 -1615 1555
rect -1648 1500 -1606 1503
rect -1658 1491 -1632 1494
rect -1608 1490 -1592 1493
rect -1592 1477 -1587 1488
rect -1519 1476 -1516 1489
rect -1500 1479 -1497 1540
rect -1412 1531 -1400 1534
rect -1488 1506 -1448 1509
rect -1447 1496 -1443 1506
rect -1500 1476 -1484 1479
rect -1364 1457 -1361 1555
rect -1342 1523 -1268 1526
rect -1342 1499 -1339 1523
rect -1320 1500 -1279 1503
rect -1281 1490 -1265 1493
rect -1264 1477 -1261 1488
rect -1192 1476 -1189 1489
rect -1173 1479 -1170 1540
rect -1085 1531 -1073 1534
rect -1161 1506 -1121 1509
rect -520 1511 -499 1514
rect -1120 1496 -1116 1506
rect -1173 1476 -1157 1479
rect -526 1456 -499 1459
rect -526 1454 -523 1456
rect -577 1451 -523 1454
rect -376 1421 -361 1424
rect -689 1399 -572 1402
rect -1618 1377 -1361 1380
rect -1746 1331 -1699 1334
rect -1618 1325 -1615 1377
rect -1648 1322 -1606 1325
rect -1658 1313 -1632 1316
rect -1608 1312 -1592 1315
rect -1592 1299 -1587 1310
rect -1519 1298 -1516 1311
rect -1500 1301 -1497 1362
rect -1412 1353 -1400 1356
rect -1488 1328 -1448 1331
rect -1447 1318 -1443 1328
rect -1500 1298 -1484 1301
rect -1729 1276 -1699 1279
rect -1364 1279 -1361 1377
rect -609 1363 -553 1366
rect -523 1363 -502 1366
rect -1342 1345 -1268 1348
rect -1342 1321 -1339 1345
rect -1320 1322 -1279 1325
rect -1281 1312 -1265 1315
rect -1264 1299 -1261 1310
rect -1192 1298 -1189 1311
rect -1173 1301 -1170 1362
rect -1085 1353 -1073 1356
rect -240 1342 -237 1440
rect -222 1384 -201 1387
rect -265 1339 -221 1342
rect -1161 1328 -1121 1331
rect -1120 1318 -1116 1328
rect -689 1323 -572 1326
rect -1173 1298 -1157 1301
rect -884 1280 -881 1318
rect -723 1297 -720 1304
rect -723 1294 -624 1297
rect -723 1288 -720 1294
rect -751 1285 -720 1288
rect -1051 1274 -917 1277
rect -751 1274 -748 1285
rect -739 1277 -699 1280
rect -627 1276 -624 1294
rect -609 1280 -553 1283
rect -810 1271 -748 1274
rect -1715 1253 -1682 1256
rect -324 1248 -321 1287
rect -265 1273 -262 1339
rect -577 1216 -507 1219
rect -329 1215 -314 1218
rect -1619 1202 -1362 1205
rect -1746 1156 -1700 1159
rect -1619 1150 -1616 1202
rect -1649 1147 -1607 1150
rect -1659 1138 -1633 1141
rect -1609 1137 -1593 1140
rect -1593 1124 -1588 1135
rect -1520 1123 -1517 1136
rect -1501 1126 -1498 1187
rect -1413 1178 -1401 1181
rect -1489 1153 -1449 1156
rect -1448 1143 -1444 1153
rect -1501 1123 -1485 1126
rect -1729 1101 -1700 1104
rect -1365 1104 -1362 1202
rect -1343 1170 -1269 1173
rect -1343 1146 -1340 1170
rect -1321 1147 -1280 1150
rect -1282 1137 -1266 1140
rect -1265 1124 -1262 1135
rect -1193 1123 -1190 1136
rect -1174 1126 -1171 1187
rect -1056 1187 -916 1190
rect -1086 1178 -1074 1181
rect -1162 1153 -1122 1156
rect -1121 1143 -1117 1153
rect -1174 1123 -1158 1126
rect -1715 1078 -1683 1081
rect -1619 1027 -1362 1030
rect -1746 981 -1700 984
rect -1619 975 -1616 1027
rect -1649 972 -1607 975
rect -1659 963 -1633 966
rect -1609 962 -1593 965
rect -1593 949 -1588 960
rect -1520 948 -1517 961
rect -1501 951 -1498 1012
rect -1413 1003 -1401 1006
rect -1489 978 -1449 981
rect -1448 968 -1444 978
rect -1501 948 -1485 951
rect -1729 926 -1700 929
rect -1365 929 -1362 1027
rect -1058 1013 -949 1016
rect -1343 995 -1269 998
rect -1343 971 -1340 995
rect -1321 972 -1280 975
rect -1282 962 -1266 965
rect -1265 949 -1262 960
rect -1193 948 -1190 961
rect -1174 951 -1171 1012
rect -1086 1003 -1074 1006
rect -1162 978 -1122 981
rect -1121 968 -1117 978
rect -1174 948 -1158 951
rect -1715 903 -1683 906
rect -1619 851 -1362 854
rect -1746 805 -1700 808
rect -1619 799 -1616 851
rect -1649 796 -1607 799
rect -1659 787 -1633 790
rect -1609 786 -1593 789
rect -1593 773 -1588 784
rect -1520 772 -1517 785
rect -1501 775 -1498 836
rect -1413 827 -1401 830
rect -1489 802 -1449 805
rect -1448 792 -1444 802
rect -1501 772 -1485 775
rect -1729 750 -1700 753
rect -1365 753 -1362 851
rect -1343 819 -1269 822
rect -1343 795 -1340 819
rect -1321 796 -1280 799
rect -1282 786 -1266 789
rect -1265 773 -1262 784
rect -1193 772 -1190 785
rect -1174 775 -1171 836
rect -1057 836 -963 839
rect -1086 827 -1074 830
rect -1162 802 -1122 805
rect -1121 792 -1117 802
rect -1174 772 -1158 775
rect -1715 727 -1683 730
rect -1619 676 -1362 679
rect -1746 630 -1717 633
rect -1729 574 -1717 577
rect -1708 512 -1705 661
rect -1619 624 -1616 676
rect -1649 621 -1607 624
rect -1659 612 -1633 615
rect -1609 611 -1593 614
rect -1593 598 -1588 609
rect -1520 597 -1517 610
rect -1501 600 -1498 661
rect -1413 652 -1401 655
rect -1489 627 -1449 630
rect -1448 617 -1444 627
rect -1501 597 -1485 600
rect -1365 578 -1362 676
rect -1343 644 -1269 647
rect -1343 620 -1340 644
rect -1321 621 -1280 624
rect -1282 611 -1266 614
rect -1265 598 -1262 609
rect -1193 597 -1190 610
rect -1174 600 -1171 661
rect -1062 661 -974 664
rect -1086 652 -1074 655
rect -1162 627 -1122 630
rect -1121 617 -1117 627
rect -1174 597 -1158 600
rect -1618 370 -1361 373
rect -1746 324 -1699 327
rect -1618 318 -1615 370
rect -1648 315 -1606 318
rect -1658 306 -1632 309
rect -1608 305 -1592 308
rect -1592 292 -1587 303
rect -1519 291 -1516 304
rect -1500 294 -1497 355
rect -1412 346 -1400 349
rect -1488 321 -1448 324
rect -1447 311 -1443 321
rect -1500 291 -1484 294
rect -1729 269 -1699 272
rect -1364 272 -1361 370
rect -1342 338 -1268 341
rect -1342 314 -1339 338
rect -1320 315 -1279 318
rect -1281 305 -1265 308
rect -1264 292 -1261 303
rect -1192 291 -1189 304
rect -1173 294 -1170 355
rect -1085 346 -1073 349
rect -1161 321 -1121 324
rect -1120 311 -1116 321
rect -1173 291 -1157 294
rect -1715 246 -1682 249
rect -1619 195 -1362 198
rect -1746 149 -1700 152
rect -1619 143 -1616 195
rect -1649 140 -1607 143
rect -1659 131 -1633 134
rect -1609 130 -1593 133
rect -1593 117 -1588 128
rect -1520 116 -1517 129
rect -1501 119 -1498 180
rect -1413 171 -1401 174
rect -1489 146 -1449 149
rect -1448 136 -1444 146
rect -1501 116 -1485 119
rect -1729 94 -1700 97
rect -1365 97 -1362 195
rect -1343 163 -1269 166
rect -1343 139 -1340 163
rect -1321 140 -1280 143
rect -1282 130 -1266 133
rect -1265 117 -1262 128
rect -1193 116 -1190 129
rect -1174 119 -1171 180
rect -1086 171 -1074 174
rect -1162 146 -1122 149
rect -1121 136 -1117 146
rect -1174 116 -1158 119
rect -1715 71 -1683 74
rect -1619 20 -1362 23
rect -1746 -26 -1700 -23
rect -1619 -32 -1616 20
rect -1649 -35 -1607 -32
rect -1659 -44 -1633 -41
rect -1609 -45 -1593 -42
rect -1593 -58 -1588 -47
rect -1520 -59 -1517 -46
rect -1501 -56 -1498 5
rect -1413 -4 -1401 -1
rect -1489 -29 -1449 -26
rect -1448 -39 -1444 -29
rect -1501 -59 -1485 -56
rect -1729 -81 -1700 -78
rect -1365 -78 -1362 20
rect -1343 -12 -1269 -9
rect -1343 -36 -1340 -12
rect -1321 -35 -1280 -32
rect -1282 -45 -1266 -42
rect -1265 -58 -1262 -47
rect -1193 -59 -1190 -46
rect -1174 -56 -1171 5
rect -1086 -4 -1074 -1
rect -1162 -29 -1122 -26
rect -1121 -39 -1117 -29
rect -1174 -59 -1158 -56
rect -1715 -104 -1683 -101
rect -1619 -156 -1362 -153
rect -1746 -202 -1700 -199
rect -1619 -208 -1616 -156
rect -1649 -211 -1607 -208
rect -1659 -220 -1633 -217
rect -1609 -221 -1593 -218
rect -1593 -234 -1588 -223
rect -1520 -235 -1517 -222
rect -1501 -232 -1498 -171
rect -1413 -180 -1401 -177
rect -1489 -205 -1449 -202
rect -1448 -215 -1444 -205
rect -1501 -235 -1485 -232
rect -1729 -257 -1700 -254
rect -1365 -254 -1362 -156
rect -1343 -188 -1269 -185
rect -1343 -212 -1340 -188
rect -1321 -211 -1280 -208
rect -1282 -221 -1266 -218
rect -1265 -234 -1262 -223
rect -1193 -235 -1190 -222
rect -1174 -232 -1171 -171
rect -1086 -180 -1074 -177
rect -1162 -205 -1122 -202
rect -1121 -215 -1117 -205
rect -1174 -235 -1158 -232
rect -1715 -280 -1683 -277
rect -1619 -331 -1362 -328
rect -1746 -377 -1717 -374
rect -1729 -433 -1717 -430
rect -1708 -495 -1705 -346
rect -1619 -383 -1616 -331
rect -1649 -386 -1607 -383
rect -1659 -395 -1633 -392
rect -1609 -396 -1593 -393
rect -1593 -409 -1588 -398
rect -1520 -410 -1517 -397
rect -1501 -407 -1498 -346
rect -1413 -355 -1401 -352
rect -1489 -380 -1449 -377
rect -1448 -390 -1444 -380
rect -1501 -410 -1485 -407
rect -1365 -429 -1362 -331
rect -1343 -363 -1269 -360
rect -1343 -387 -1340 -363
rect -1321 -386 -1280 -383
rect -1282 -396 -1266 -393
rect -1265 -409 -1262 -398
rect -1193 -410 -1190 -397
rect -1174 -407 -1171 -346
rect -1086 -355 -1074 -352
rect -1162 -380 -1122 -377
rect -1121 -390 -1117 -380
rect -1174 -410 -1158 -407
rect -977 -407 -974 661
rect -966 95 -963 836
rect -952 542 -949 1013
rect -932 909 -929 1187
rect -240 1172 -237 1339
rect -157 1341 -154 1379
rect 4 1358 7 1365
rect 4 1355 103 1358
rect 4 1349 7 1355
rect -24 1346 7 1349
rect -24 1335 -21 1346
rect -12 1338 28 1341
rect 100 1337 103 1355
rect -83 1332 -21 1335
rect -201 1289 -180 1292
rect -191 1253 -188 1275
rect -191 1250 -70 1253
rect -129 1174 -126 1212
rect -577 1161 -505 1164
rect -389 1160 -353 1163
rect -541 1148 -493 1151
rect -693 1033 -572 1036
rect -609 997 -553 1000
rect -693 957 -572 960
rect -888 914 -885 952
rect -727 931 -724 938
rect -541 940 -538 1148
rect -356 1085 -353 1160
rect -341 1138 -338 1158
rect -411 1082 -353 1085
rect -356 1055 -353 1082
rect -368 1051 -357 1054
rect -368 1017 -365 1051
rect -152 1017 -149 1119
rect -368 1014 -149 1017
rect -523 997 -467 1000
rect -116 990 -113 1139
rect -154 986 -117 989
rect -92 979 -89 1190
rect -476 976 -89 979
rect -541 937 -499 940
rect -727 928 -628 931
rect -727 922 -724 928
rect -755 919 -724 922
rect -755 908 -752 919
rect -743 911 -703 914
rect -631 910 -628 928
rect -609 914 -553 917
rect -814 905 -752 908
rect -539 852 -536 900
rect -502 824 -499 937
rect -476 857 -473 976
rect -73 968 -70 1250
rect 32 1191 35 1198
rect 32 1188 131 1191
rect 32 1182 35 1188
rect 4 1179 35 1182
rect 4 1168 7 1179
rect 16 1171 56 1174
rect 128 1170 131 1188
rect -55 1165 7 1168
rect -468 965 -70 968
rect -468 841 -465 965
rect -64 894 -61 914
rect -315 861 -249 864
rect -21 855 -18 893
rect 140 872 143 879
rect 140 869 239 872
rect 140 863 143 869
rect 112 860 143 863
rect 112 849 115 860
rect 124 852 164 855
rect 236 851 239 869
rect 53 846 115 849
rect -333 826 -280 829
rect -577 806 -467 809
rect -339 806 -233 809
rect -502 776 -499 786
rect -502 773 -475 776
rect -497 765 -479 768
rect -343 739 -340 805
rect -236 803 -127 806
rect -53 799 -50 815
rect -328 757 -293 760
rect -347 736 -340 739
rect -693 675 -572 678
rect -474 645 -471 684
rect -343 661 -340 736
rect -314 681 -285 684
rect -369 658 -340 661
rect -609 639 -553 642
rect -535 626 -480 629
rect -693 599 -572 602
rect -888 556 -885 594
rect -727 573 -724 580
rect -727 570 -628 573
rect -727 564 -724 570
rect -755 561 -724 564
rect -755 550 -752 561
rect -743 553 -703 556
rect -631 552 -628 570
rect -609 556 -553 559
rect -814 547 -752 550
rect -693 228 -572 231
rect -609 192 -553 195
rect -693 152 -572 155
rect -888 109 -885 147
rect -727 126 -724 133
rect -727 123 -628 126
rect -727 117 -724 123
rect -755 114 -724 117
rect -755 103 -752 114
rect -743 106 -703 109
rect -631 105 -628 123
rect -609 109 -553 112
rect -814 100 -752 103
rect -693 -275 -572 -272
rect -609 -311 -553 -308
rect -693 -351 -572 -348
rect -888 -394 -885 -356
rect -727 -377 -724 -370
rect -727 -380 -628 -377
rect -727 -386 -724 -380
rect -755 -389 -724 -386
rect -755 -400 -752 -389
rect -743 -397 -703 -394
rect -631 -398 -628 -380
rect -609 -394 -553 -391
rect -814 -403 -752 -400
<< labels >>
rlabel metal1 -1771 1322 -1751 1343 7 A0
rlabel metal1 -1771 1147 -1751 1168 7 A1
rlabel metal1 -1771 972 -1751 993 7 A2
rlabel metal1 -1771 796 -1751 817 7 A3
rlabel metal1 -1771 621 -1751 642 7 A4
rlabel metal1 -1737 -518 -1734 -515 2 CLK
rlabel metal1 -1708 -518 -1705 -515 1 VDD
rlabel metal1 -1723 -518 -1720 -515 2 GND
rlabel metal1 -1771 315 -1751 336 7 B0
rlabel metal1 -1771 140 -1751 161 7 B1
rlabel metal1 -1771 -35 -1751 -14 7 B2
rlabel metal1 -1771 -211 -1751 -190 7 B3
rlabel metal1 -1771 -386 -1751 -365 7 B4
rlabel metal1 -548 -402 -528 -381 7 P4
rlabel metal1 -548 -319 -528 -298 7 G4
rlabel metal1 -548 101 -528 122 7 P3
rlabel metal1 -548 184 -528 205 7 G3
rlabel metal1 -548 547 -528 568 7 P2
rlabel metal1 -548 630 -528 651 7 G2
rlabel metal1 -548 905 -528 926 7 P1
rlabel metal1 -548 989 -528 1010 7 G1
rlabel metal1 -548 1271 -528 1292 7 P0
rlabel metal1 -548 1354 -528 1375 7 G0
rlabel metal1 -1751 1500 -1731 1521 1 Cin
rlabel metal1 117 1332 137 1353 1 S0
rlabel metal1 -176 1066 -172 1070 1 C1
rlabel metal1 141 1165 161 1186 1 S1
rlabel metal1 -90 823 -86 827 1 C2
rlabel metal1 249 846 269 867 1 S2
<< end >>
