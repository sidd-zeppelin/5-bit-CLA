* NGSPICE file created from NOR6.ext - technology: scmos

.global Vdd Gnd 


* Top level circuit NOR6

M1000 GND B OUT Gnd cmosn w=0.9u l=0.18u
+  ad=1.782p pd=11.16u as=1.458p ps=8.64u
M1001 a_19_n4# A VDD Vdd cmosp w=10.8u l=0.18u
+  ad=5.832p pd=22.68u as=4.86p ps=22.5u
M1002 GND D OUT Gnd cmosn w=0.9u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1003 a_19_28# E a_19_20# Vdd cmosp w=10.8u l=0.18u
+  ad=5.832p pd=22.68u as=5.832p ps=22.68u
M1004 a_19_4# B a_19_n4# Vdd cmosp w=10.8u l=0.18u
+  ad=5.832p pd=22.68u as=0p ps=0u
M1005 OUT A GND Gnd cmosn w=0.9u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1006 a_19_12# C a_19_4# Vdd cmosp w=10.8u l=0.18u
+  ad=5.832p pd=22.68u as=0p ps=0u
M1007 OUT E GND Gnd cmosn w=0.9u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1008 OUT F a_19_28# Vdd cmosp w=10.8u l=0.18u
+  ad=4.86p pd=22.5u as=0p ps=0u
M1009 OUT C GND Gnd cmosn w=0.9u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1010 GND F OUT Gnd cmosn w=0.9u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_19_20# D a_19_12# Vdd cmosp w=10.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
.end

