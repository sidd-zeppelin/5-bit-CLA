* SPICE3 file created from NAND2.ext - technology: scmos

.option scale=0.09u

M1000 OUT A VDD w_n6_26# cmosp w=20 l=2
+  ad=120 pd=52 as=200 ps=100
M1001 VDD B OUT w_n6_26# cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1002 OUT B a_7_n1# Gnd cmosn w=20 l=2
+  ad=100 pd=50 as=120 ps=52
M1003 a_7_n1# A GND Gnd cmosn w=20 l=2
+  ad=0 pd=0 as=100 ps=50
