* SPICE3 file created from NOR5.ext - technology: scmos

.option scale=0.09u

M1000 a_31_22# D a_23_22# w_n6_16# cmosp w=100 l=2
+  ad=600 pd=212 as=600 ps=212
M1001 a_7_22# A VDD w_n6_16# cmosp w=100 l=2
+  ad=600 pd=212 as=500 ps=210
M1002 GND D OUT Gnd cmosn w=10 l=2
+  ad=170 pd=94 as=170 ps=94
M1003 GND B OUT Gnd cmosn w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 a_15_22# B a_7_22# w_n6_16# cmosp w=100 l=2
+  ad=600 pd=212 as=0 ps=0
M1005 OUT A GND Gnd cmosn w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 OUT E GND Gnd cmosn w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1007 OUT E a_31_22# w_n6_16# cmosp w=100 l=2
+  ad=500 pd=210 as=0 ps=0
M1008 OUT C GND Gnd cmosn w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1009 a_23_22# C a_15_22# w_n6_16# cmosp w=100 l=2
+  ad=0 pd=0 as=0 ps=0
C0 w_n6_16# Gnd 6.30fF
