* SPICE3 file created from AND4.ext - technology: scmos

.option scale=0.09u

M1000 a_49_21# B a_49_13# Gnd cmosn w=40 l=2
+  ad=240 pd=92 as=240 ps=92
M1001 VDD B a_17_13# w_11_0# cmosp w=20 l=2
+  ad=420 pd=202 as=240 ps=104
M1002 a_49_29# C a_49_21# Gnd cmosn w=40 l=2
+  ad=240 pd=92 as=0 ps=0
M1003 a_17_13# C VDD w_11_0# cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 a_49_13# A GND Gnd cmosn w=40 l=2
+  ad=0 pd=0 as=250 ps=120
M1005 a_17_13# A VDD w_11_0# cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 OUT a_17_13# VDD w_103_23# cmosp w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1007 a_17_13# D a_49_29# Gnd cmosn w=40 l=2
+  ad=200 pd=90 as=0 ps=0
M1008 VDD D a_17_13# w_11_0# cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1009 OUT a_17_13# GND Gnd cmosn w=10 l=2
+  ad=50 pd=30 as=0 ps=0
