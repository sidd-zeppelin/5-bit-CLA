magic
tech scmos
timestamp 1763744018
<< nwell >>
rect 11 0 83 40
rect 113 19 137 51
<< ntransistor >>
rect 89 27 99 29
rect 89 19 99 21
rect 89 11 99 13
rect 124 -1 126 9
<< ptransistor >>
rect 17 27 77 29
rect 124 25 126 45
rect 17 19 77 21
rect 17 11 77 13
<< ndiffusion >>
rect 89 29 99 30
rect 89 26 99 27
rect 89 21 99 22
rect 89 18 99 19
rect 89 13 99 14
rect 89 10 99 11
rect 123 -1 124 9
rect 126 -1 127 9
<< pdiffusion >>
rect 17 29 77 30
rect 17 26 77 27
rect 17 21 77 22
rect 123 25 124 45
rect 126 25 127 45
rect 17 18 77 19
rect 17 13 77 14
rect 17 10 77 11
<< ndcontact >>
rect 89 30 99 34
rect 89 22 99 26
rect 89 14 99 18
rect 89 6 99 10
rect 119 -1 123 9
rect 127 -1 131 9
<< pdcontact >>
rect 17 30 77 34
rect 17 22 77 26
rect 119 25 123 45
rect 127 25 131 45
rect 17 14 77 18
rect 17 6 77 10
<< polysilicon >>
rect 124 45 126 48
rect 8 27 17 29
rect 77 27 89 29
rect 99 27 102 29
rect 8 19 17 21
rect 77 19 89 21
rect 99 19 102 21
rect 8 11 17 13
rect 77 11 89 13
rect 99 11 102 13
rect 124 9 126 25
rect 124 -4 126 -1
<< polycontact >>
rect 4 26 8 30
rect 4 18 8 22
rect 4 10 8 14
rect 120 12 124 16
<< metal1 >>
rect 0 48 137 51
rect 0 26 4 30
rect 0 18 4 22
rect 0 10 4 14
rect 11 10 14 48
rect 119 45 123 48
rect 83 37 113 40
rect 83 34 86 37
rect 77 30 89 34
rect 83 18 86 30
rect 102 26 105 34
rect 99 22 105 26
rect 83 14 89 18
rect 102 10 105 22
rect 110 16 113 37
rect 127 16 131 25
rect 110 12 120 16
rect 127 12 137 16
rect 11 6 17 10
rect 99 6 105 10
rect 127 9 131 12
rect 11 0 14 6
rect 102 -4 105 6
rect 119 -4 123 -1
rect 0 -7 131 -4
<< labels >>
rlabel metal1 0 10 4 14 3 A
rlabel metal1 0 18 4 22 3 B
rlabel metal1 0 26 4 30 3 C
rlabel metal1 133 12 137 16 7 OUT
rlabel metal1 0 48 3 51 4 VDD
rlabel metal1 0 -7 3 -4 2 GND
<< end >>
