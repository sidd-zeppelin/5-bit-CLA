* SPICE3 file created from AND2.ext - technology: scmos

.option scale=0.09u

M1000 OUT a_n21_n16# VDD w_46_n8# cmosp w=20 l=2
+  ad=100 pd=50 as=300 ps=150
M1001 a_n21_n16# A VDD w_n27_n29# cmosp w=20 l=2
+  ad=120 pd=52 as=0 ps=0
M1002 VDD B a_n21_n16# w_n27_n29# cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 a_12_n16# A GND Gnd cmosn w=20 l=2
+  ad=120 pd=52 as=150 ps=80
M1004 OUT a_n21_n16# GND Gnd cmosn w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1005 a_n21_n16# B a_12_n16# Gnd cmosn w=20 l=2
+  ad=100 pd=50 as=0 ps=0
