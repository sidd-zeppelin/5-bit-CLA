magic
tech scmos
timestamp 1764774576
<< nwell >>
rect 649 1271 681 1303
rect 714 1271 746 1303
rect 791 1271 823 1303
rect 856 1271 888 1303
rect 931 1271 963 1303
rect 996 1271 1028 1303
rect 1076 1271 1108 1303
rect 1141 1271 1173 1303
rect 1221 1271 1253 1303
rect 1286 1271 1318 1303
rect 1366 1271 1398 1303
rect 1431 1271 1463 1303
rect 667 1165 699 1197
rect 714 1165 746 1197
rect 809 1165 841 1197
rect 856 1165 888 1197
rect 949 1165 981 1197
rect 996 1165 1028 1197
rect 1094 1165 1126 1197
rect 1141 1165 1173 1197
rect 1239 1165 1271 1197
rect 1286 1165 1318 1197
rect 1384 1165 1416 1197
rect 1431 1165 1463 1197
rect -580 1090 -548 1122
rect -474 1108 -442 1140
rect -253 1090 -221 1122
rect -147 1108 -115 1140
rect 699 1120 731 1144
rect 841 1120 873 1144
rect 981 1120 1013 1144
rect 1126 1120 1158 1144
rect 1271 1120 1303 1144
rect 1416 1120 1448 1144
rect -676 1058 -652 1090
rect -625 1058 -601 1090
rect -580 1043 -548 1075
rect -474 1043 -442 1075
rect -348 1058 -324 1090
rect -298 1058 -274 1090
rect -253 1043 -221 1075
rect -147 1043 -115 1075
rect 699 1070 731 1094
rect 841 1070 873 1094
rect 981 1070 1013 1094
rect 1126 1070 1158 1094
rect 1271 1070 1303 1094
rect 1416 1070 1448 1094
rect 410 1006 442 1038
rect -1240 930 -1208 962
rect -1134 948 -1102 980
rect -913 930 -881 962
rect -807 948 -775 980
rect -1336 898 -1312 930
rect -1285 898 -1261 930
rect -1240 883 -1208 915
rect -1134 883 -1102 915
rect -1008 898 -984 930
rect -958 898 -934 930
rect -581 926 -549 958
rect -475 944 -443 976
rect -254 926 -222 958
rect -148 944 -116 976
rect 319 972 351 1004
rect 410 950 442 982
rect 506 972 538 1004
rect -913 883 -881 915
rect -807 883 -775 915
rect -677 894 -653 926
rect -626 894 -602 926
rect -581 879 -549 911
rect -475 879 -443 911
rect -349 894 -325 926
rect -299 894 -275 926
rect 159 918 191 950
rect 649 944 681 976
rect 714 944 746 976
rect 791 944 823 976
rect 856 944 888 976
rect 931 944 963 976
rect 996 944 1028 976
rect 1076 944 1108 976
rect 1141 944 1173 976
rect 1221 944 1253 976
rect 1286 944 1318 976
rect 1366 944 1398 976
rect 1431 944 1463 976
rect -254 879 -222 911
rect -148 879 -116 911
rect 68 884 100 916
rect 159 862 191 894
rect 255 884 287 916
rect 362 865 394 897
rect 435 886 459 918
rect 480 864 532 896
rect 563 886 587 918
rect 53 804 85 836
rect 126 825 150 857
rect 667 838 699 870
rect 714 838 746 870
rect 809 838 841 870
rect 856 838 888 870
rect 949 838 981 870
rect 996 838 1028 870
rect 1094 838 1126 870
rect 1141 838 1173 870
rect 1239 838 1271 870
rect 1286 838 1318 870
rect 1384 838 1416 870
rect 1431 838 1463 870
rect 285 779 317 811
rect 358 800 382 832
rect 409 774 481 814
rect 511 793 535 825
rect 699 793 731 817
rect 841 793 873 817
rect 981 793 1013 817
rect 1126 793 1158 817
rect 1271 793 1303 817
rect 1416 793 1448 817
rect -1240 691 -1208 723
rect -1134 709 -1102 741
rect -913 691 -881 723
rect -807 709 -775 741
rect -1336 659 -1312 691
rect -1285 659 -1261 691
rect -1240 644 -1208 676
rect -1134 644 -1102 676
rect -1008 659 -984 691
rect -958 659 -934 691
rect -581 690 -549 722
rect -475 708 -443 740
rect -254 690 -222 722
rect -148 708 -116 740
rect 158 738 190 770
rect 699 742 731 766
rect 841 742 873 766
rect 981 742 1013 766
rect 1126 742 1158 766
rect 1271 742 1303 766
rect 1416 742 1448 766
rect 67 704 99 736
rect -913 644 -881 676
rect -807 644 -775 676
rect -677 658 -653 690
rect -626 658 -602 690
rect -581 643 -549 675
rect -475 643 -443 675
rect -349 658 -325 690
rect -299 658 -275 690
rect 158 682 190 714
rect 254 704 286 736
rect 368 689 400 729
rect 450 707 474 739
rect -254 643 -222 675
rect -148 643 -116 675
rect 52 624 84 656
rect 125 645 149 677
rect 649 651 681 683
rect 290 611 322 643
rect 558 617 590 649
rect 199 577 231 609
rect 290 555 322 587
rect 386 577 418 609
rect 649 595 681 627
rect 745 617 777 649
rect -1240 477 -1208 509
rect -1134 495 -1102 527
rect -913 477 -881 509
rect -807 495 -775 527
rect -1336 445 -1312 477
rect -1285 445 -1261 477
rect -1240 430 -1208 462
rect -1134 430 -1102 462
rect -1008 445 -984 477
rect -958 445 -934 477
rect -581 476 -549 508
rect -475 494 -443 526
rect -254 476 -222 508
rect -148 494 -116 526
rect 158 484 190 516
rect 542 513 574 545
rect 615 534 639 566
rect -913 430 -881 462
rect -807 430 -775 462
rect -677 444 -653 476
rect -626 444 -602 476
rect -581 429 -549 461
rect -475 429 -443 461
rect -349 444 -325 476
rect -299 444 -275 476
rect -254 429 -222 461
rect -148 429 -116 461
rect 67 450 99 482
rect 158 428 190 460
rect 254 450 286 482
rect 373 446 405 494
rect 465 469 489 501
rect 542 452 574 492
rect 624 470 648 502
rect 689 460 781 508
rect 812 481 836 513
rect 52 370 84 402
rect 125 391 149 423
rect 719 392 751 424
rect 792 413 816 445
rect 159 302 191 334
rect 301 325 333 381
rect 379 357 403 389
rect 437 335 469 383
rect 529 358 553 390
rect 583 340 615 380
rect 665 358 689 390
rect 729 304 841 360
rect 870 337 894 369
rect -1240 238 -1208 270
rect -1134 256 -1102 288
rect -913 238 -881 270
rect -807 256 -775 288
rect -1336 206 -1312 238
rect -1285 206 -1261 238
rect -1240 191 -1208 223
rect -1134 191 -1102 223
rect -1008 206 -984 238
rect -958 206 -934 238
rect -581 237 -549 269
rect -475 255 -443 287
rect -254 237 -222 269
rect -148 255 -116 287
rect 68 268 100 300
rect 159 246 191 278
rect 255 268 287 300
rect -913 191 -881 223
rect -807 191 -775 223
rect -677 205 -653 237
rect -626 205 -602 237
rect -581 190 -549 222
rect -475 190 -443 222
rect -349 205 -325 237
rect -299 205 -275 237
rect -254 190 -222 222
rect -148 190 -116 222
rect 53 188 85 220
rect 126 209 150 241
rect 482 233 514 265
rect 391 199 423 231
rect 482 177 514 209
rect 578 199 610 231
rect 700 172 732 212
rect 782 190 806 222
rect 846 192 878 224
rect 919 213 943 245
rect 1107 230 1139 262
rect 1016 196 1048 228
rect 1107 174 1139 206
rect 1203 196 1235 228
rect 160 119 192 151
rect -1240 51 -1208 83
rect -1134 69 -1102 101
rect -913 51 -881 83
rect -807 69 -775 101
rect -1336 19 -1312 51
rect -1285 19 -1261 51
rect -1240 4 -1208 36
rect -1134 4 -1102 36
rect -1008 19 -984 51
rect -958 19 -934 51
rect -581 50 -549 82
rect -475 68 -443 100
rect -254 50 -222 82
rect -148 68 -116 100
rect 69 85 101 117
rect 160 63 192 95
rect 256 85 288 117
rect 382 77 405 141
rect 464 110 488 142
rect 519 87 551 143
rect 597 119 621 151
rect 647 87 679 135
rect 739 110 763 142
rect 858 75 990 139
rect 1028 108 1052 140
rect -913 4 -881 36
rect -807 4 -775 36
rect -677 18 -653 50
rect -626 18 -602 50
rect -581 3 -549 35
rect -475 3 -443 35
rect -349 18 -325 50
rect -299 18 -275 50
rect -254 3 -222 35
rect -148 3 -116 35
rect 54 5 86 37
rect 127 26 151 58
<< polysilicon >>
rect 660 1333 662 1336
rect 668 1333 670 1336
rect 725 1333 727 1336
rect 733 1333 735 1336
rect 802 1333 804 1336
rect 810 1333 812 1336
rect 867 1333 869 1336
rect 875 1333 877 1336
rect 942 1333 944 1336
rect 950 1333 952 1336
rect 1007 1333 1009 1336
rect 1015 1333 1017 1336
rect 1087 1333 1089 1336
rect 1095 1333 1097 1336
rect 1152 1333 1154 1336
rect 1160 1333 1162 1336
rect 1232 1333 1234 1336
rect 1240 1333 1242 1336
rect 1297 1333 1299 1336
rect 1305 1333 1307 1336
rect 1377 1333 1379 1336
rect 1385 1333 1387 1336
rect 1442 1333 1444 1336
rect 1450 1333 1452 1336
rect 660 1297 662 1313
rect 668 1297 670 1313
rect 725 1297 727 1313
rect 733 1297 735 1313
rect 802 1297 804 1313
rect 810 1297 812 1313
rect 867 1297 869 1313
rect 875 1297 877 1313
rect 942 1297 944 1313
rect 950 1297 952 1313
rect 1007 1297 1009 1313
rect 1015 1297 1017 1313
rect 1087 1297 1089 1313
rect 1095 1297 1097 1313
rect 1152 1297 1154 1313
rect 1160 1297 1162 1313
rect 1232 1297 1234 1313
rect 1240 1297 1242 1313
rect 1297 1297 1299 1313
rect 1305 1297 1307 1313
rect 1377 1297 1379 1313
rect 1385 1297 1387 1313
rect 1442 1297 1444 1313
rect 1450 1297 1452 1313
rect 660 1265 662 1277
rect 668 1265 670 1277
rect 725 1265 727 1277
rect 733 1265 735 1277
rect 802 1265 804 1277
rect 810 1265 812 1277
rect 867 1265 869 1277
rect 875 1265 877 1277
rect 942 1265 944 1277
rect 950 1265 952 1277
rect 1007 1265 1009 1277
rect 1015 1265 1017 1277
rect 1087 1265 1089 1277
rect 1095 1265 1097 1277
rect 1152 1265 1154 1277
rect 1160 1265 1162 1277
rect 1232 1265 1234 1277
rect 1240 1265 1242 1277
rect 1297 1265 1299 1277
rect 1305 1265 1307 1277
rect 1377 1265 1379 1277
rect 1385 1265 1387 1277
rect 1442 1265 1444 1277
rect 1450 1265 1452 1277
rect 678 1227 680 1230
rect 686 1227 688 1230
rect 725 1227 727 1230
rect 733 1227 735 1230
rect 820 1227 822 1230
rect 828 1227 830 1230
rect 867 1227 869 1230
rect 875 1227 877 1230
rect 960 1227 962 1230
rect 968 1227 970 1230
rect 1007 1227 1009 1230
rect 1015 1227 1017 1230
rect 1105 1227 1107 1230
rect 1113 1227 1115 1230
rect 1152 1227 1154 1230
rect 1160 1227 1162 1230
rect 1250 1227 1252 1230
rect 1258 1227 1260 1230
rect 1297 1227 1299 1230
rect 1305 1227 1307 1230
rect 1395 1227 1397 1230
rect 1403 1227 1405 1230
rect 1442 1227 1444 1230
rect 1450 1227 1452 1230
rect 678 1191 680 1207
rect 686 1191 688 1207
rect 725 1191 727 1207
rect 733 1191 735 1207
rect 820 1191 822 1207
rect 828 1191 830 1207
rect 867 1191 869 1207
rect 875 1191 877 1207
rect 960 1191 962 1207
rect 968 1191 970 1207
rect 1007 1191 1009 1207
rect 1015 1191 1017 1207
rect 1105 1191 1107 1207
rect 1113 1191 1115 1207
rect 1152 1191 1154 1207
rect 1160 1191 1162 1207
rect 1250 1191 1252 1207
rect 1258 1191 1260 1207
rect 1297 1191 1299 1207
rect 1305 1191 1307 1207
rect 1395 1191 1397 1207
rect 1403 1191 1405 1207
rect 1442 1191 1444 1207
rect 1450 1191 1452 1207
rect 678 1159 680 1171
rect 686 1159 688 1171
rect 725 1159 727 1171
rect 733 1159 735 1171
rect 820 1159 822 1171
rect 828 1159 830 1171
rect 867 1159 869 1171
rect 875 1159 877 1171
rect 960 1159 962 1171
rect 968 1159 970 1171
rect 1007 1159 1009 1171
rect 1015 1159 1017 1171
rect 1105 1159 1107 1171
rect 1113 1159 1115 1171
rect 1152 1159 1154 1171
rect 1160 1159 1162 1171
rect 1250 1159 1252 1171
rect 1258 1159 1260 1171
rect 1297 1159 1299 1171
rect 1305 1159 1307 1171
rect 1395 1159 1397 1171
rect 1403 1159 1405 1171
rect 1442 1159 1444 1171
rect 1450 1159 1452 1171
rect -480 1127 -468 1129
rect -448 1127 -432 1129
rect -412 1127 -409 1129
rect 702 1131 705 1133
rect 725 1131 739 1133
rect 749 1131 752 1133
rect 844 1131 847 1133
rect 867 1131 881 1133
rect 891 1131 894 1133
rect 984 1131 987 1133
rect 1007 1131 1021 1133
rect 1031 1131 1034 1133
rect 1129 1131 1132 1133
rect 1152 1131 1166 1133
rect 1176 1131 1179 1133
rect 1274 1131 1277 1133
rect 1297 1131 1311 1133
rect 1321 1131 1324 1133
rect 1419 1131 1422 1133
rect 1442 1131 1456 1133
rect 1466 1131 1469 1133
rect -153 1127 -141 1129
rect -121 1127 -105 1129
rect -85 1127 -82 1129
rect -480 1119 -468 1121
rect -448 1119 -432 1121
rect -412 1119 -409 1121
rect -153 1119 -141 1121
rect -121 1119 -105 1121
rect -85 1119 -82 1121
rect -586 1109 -574 1111
rect -554 1109 -538 1111
rect -518 1109 -515 1111
rect -259 1109 -247 1111
rect -227 1109 -211 1111
rect -191 1109 -188 1111
rect -586 1101 -574 1103
rect -554 1101 -538 1103
rect -518 1101 -515 1103
rect -259 1101 -247 1103
rect -227 1101 -211 1103
rect -191 1101 -188 1103
rect -665 1084 -663 1087
rect -614 1084 -612 1087
rect -337 1084 -335 1087
rect -287 1084 -285 1087
rect -665 1050 -663 1064
rect -614 1050 -612 1064
rect -586 1062 -574 1064
rect -554 1062 -538 1064
rect -518 1062 -515 1064
rect 702 1081 705 1083
rect 725 1081 739 1083
rect 749 1081 752 1083
rect 844 1081 847 1083
rect 867 1081 881 1083
rect 891 1081 894 1083
rect 984 1081 987 1083
rect 1007 1081 1021 1083
rect 1031 1081 1034 1083
rect 1129 1081 1132 1083
rect 1152 1081 1166 1083
rect 1176 1081 1179 1083
rect 1274 1081 1277 1083
rect 1297 1081 1311 1083
rect 1321 1081 1324 1083
rect 1419 1081 1422 1083
rect 1442 1081 1456 1083
rect 1466 1081 1469 1083
rect -480 1062 -468 1064
rect -448 1062 -432 1064
rect -412 1062 -409 1064
rect -586 1054 -574 1056
rect -554 1054 -538 1056
rect -518 1054 -515 1056
rect -480 1054 -468 1056
rect -448 1054 -432 1056
rect -412 1054 -409 1056
rect -337 1050 -335 1064
rect -287 1050 -285 1064
rect -259 1062 -247 1064
rect -227 1062 -211 1064
rect -191 1062 -188 1064
rect -153 1062 -141 1064
rect -121 1062 -105 1064
rect -85 1062 -82 1064
rect -259 1054 -247 1056
rect -227 1054 -211 1056
rect -191 1054 -188 1056
rect -153 1054 -141 1056
rect -121 1054 -105 1056
rect -85 1054 -82 1056
rect -665 1037 -663 1040
rect -614 1037 -612 1040
rect -337 1037 -335 1040
rect -287 1037 -285 1040
rect 404 1025 416 1027
rect 436 1025 452 1027
rect 472 1025 475 1027
rect 404 1017 416 1019
rect 436 1017 452 1019
rect 472 1017 475 1019
rect 660 1006 662 1009
rect 668 1006 670 1009
rect 725 1006 727 1009
rect 733 1006 735 1009
rect 802 1006 804 1009
rect 810 1006 812 1009
rect 867 1006 869 1009
rect 875 1006 877 1009
rect 942 1006 944 1009
rect 950 1006 952 1009
rect 1007 1006 1009 1009
rect 1015 1006 1017 1009
rect 1087 1006 1089 1009
rect 1095 1006 1097 1009
rect 1152 1006 1154 1009
rect 1160 1006 1162 1009
rect 1232 1006 1234 1009
rect 1240 1006 1242 1009
rect 1297 1006 1299 1009
rect 1305 1006 1307 1009
rect 1377 1006 1379 1009
rect 1385 1006 1387 1009
rect 1442 1006 1444 1009
rect 1450 1006 1452 1009
rect 313 991 325 993
rect 345 991 361 993
rect 381 991 384 993
rect 500 991 512 993
rect 532 991 548 993
rect 568 991 571 993
rect 313 983 325 985
rect 345 983 361 985
rect 381 983 384 985
rect 500 983 512 985
rect 532 983 548 985
rect 568 983 571 985
rect -1140 967 -1128 969
rect -1108 967 -1092 969
rect -1072 967 -1069 969
rect -813 967 -801 969
rect -781 967 -765 969
rect -745 967 -742 969
rect -1140 959 -1128 961
rect -1108 959 -1092 961
rect -1072 959 -1069 961
rect -481 963 -469 965
rect -449 963 -433 965
rect -413 963 -410 965
rect -813 959 -801 961
rect -781 959 -765 961
rect -745 959 -742 961
rect -1246 949 -1234 951
rect -1214 949 -1198 951
rect -1178 949 -1175 951
rect 404 969 416 971
rect 436 969 452 971
rect 472 969 475 971
rect 660 970 662 986
rect 668 970 670 986
rect 725 970 727 986
rect 733 970 735 986
rect 802 970 804 986
rect 810 970 812 986
rect 867 970 869 986
rect 875 970 877 986
rect 942 970 944 986
rect 950 970 952 986
rect 1007 970 1009 986
rect 1015 970 1017 986
rect 1087 970 1089 986
rect 1095 970 1097 986
rect 1152 970 1154 986
rect 1160 970 1162 986
rect 1232 970 1234 986
rect 1240 970 1242 986
rect 1297 970 1299 986
rect 1305 970 1307 986
rect 1377 970 1379 986
rect 1385 970 1387 986
rect 1442 970 1444 986
rect 1450 970 1452 986
rect -154 963 -142 965
rect -122 963 -106 965
rect -86 963 -83 965
rect -481 955 -469 957
rect -449 955 -433 957
rect -413 955 -410 957
rect -919 949 -907 951
rect -887 949 -871 951
rect -851 949 -848 951
rect -1246 941 -1234 943
rect -1214 941 -1198 943
rect -1178 941 -1175 943
rect 404 961 416 963
rect 436 961 452 963
rect 472 961 475 963
rect -154 955 -142 957
rect -122 955 -106 957
rect -86 955 -83 957
rect -587 945 -575 947
rect -555 945 -539 947
rect -519 945 -516 947
rect -919 941 -907 943
rect -887 941 -871 943
rect -851 941 -848 943
rect -260 945 -248 947
rect -228 945 -212 947
rect -192 945 -189 947
rect -587 937 -575 939
rect -555 937 -539 939
rect -519 937 -516 939
rect -260 937 -248 939
rect -228 937 -212 939
rect -192 937 -189 939
rect 153 937 165 939
rect 185 937 201 939
rect 221 937 224 939
rect 660 938 662 950
rect 668 938 670 950
rect 725 938 727 950
rect 733 938 735 950
rect 802 938 804 950
rect 810 938 812 950
rect 867 938 869 950
rect 875 938 877 950
rect 942 938 944 950
rect 950 938 952 950
rect 1007 938 1009 950
rect 1015 938 1017 950
rect 1087 938 1089 950
rect 1095 938 1097 950
rect 1152 938 1154 950
rect 1160 938 1162 950
rect 1232 938 1234 950
rect 1240 938 1242 950
rect 1297 938 1299 950
rect 1305 938 1307 950
rect 1377 938 1379 950
rect 1385 938 1387 950
rect 1442 938 1444 950
rect 1450 938 1452 950
rect 153 929 165 931
rect 185 929 201 931
rect 221 929 224 931
rect -1325 924 -1323 927
rect -1274 924 -1272 927
rect -997 924 -995 927
rect -947 924 -945 927
rect -1325 890 -1323 904
rect -1274 890 -1272 904
rect -1246 902 -1234 904
rect -1214 902 -1198 904
rect -1178 902 -1175 904
rect -666 920 -664 923
rect -615 920 -613 923
rect -338 920 -336 923
rect -288 920 -286 923
rect -1140 902 -1128 904
rect -1108 902 -1092 904
rect -1072 902 -1069 904
rect -1246 894 -1234 896
rect -1214 894 -1198 896
rect -1178 894 -1175 896
rect -1140 894 -1128 896
rect -1108 894 -1092 896
rect -1072 894 -1069 896
rect -997 890 -995 904
rect -947 890 -945 904
rect -919 902 -907 904
rect -887 902 -871 904
rect -851 902 -848 904
rect -813 902 -801 904
rect -781 902 -765 904
rect -745 902 -742 904
rect -919 894 -907 896
rect -887 894 -871 896
rect -851 894 -848 896
rect -813 894 -801 896
rect -781 894 -765 896
rect -745 894 -742 896
rect -666 886 -664 900
rect -615 886 -613 900
rect -587 898 -575 900
rect -555 898 -539 900
rect -519 898 -516 900
rect 446 912 448 915
rect 574 912 576 915
rect -481 898 -469 900
rect -449 898 -433 900
rect -413 898 -410 900
rect -587 890 -575 892
rect -555 890 -539 892
rect -519 890 -516 892
rect -1325 877 -1323 880
rect -1274 877 -1272 880
rect -997 877 -995 880
rect -947 877 -945 880
rect -481 890 -469 892
rect -449 890 -433 892
rect -413 890 -410 892
rect -338 886 -336 900
rect -288 886 -286 900
rect -260 898 -248 900
rect -228 898 -212 900
rect -192 898 -189 900
rect 62 903 74 905
rect 94 903 110 905
rect 130 903 133 905
rect -154 898 -142 900
rect -122 898 -106 900
rect -86 898 -83 900
rect -260 890 -248 892
rect -228 890 -212 892
rect -192 890 -189 892
rect 249 903 261 905
rect 281 903 297 905
rect 317 903 320 905
rect 62 895 74 897
rect 94 895 110 897
rect 130 895 133 897
rect -154 890 -142 892
rect -122 890 -106 892
rect -86 890 -83 892
rect 249 895 261 897
rect 281 895 297 897
rect 317 895 320 897
rect 678 900 680 903
rect 686 900 688 903
rect 725 900 727 903
rect 733 900 735 903
rect 820 900 822 903
rect 828 900 830 903
rect 867 900 869 903
rect 875 900 877 903
rect 960 900 962 903
rect 968 900 970 903
rect 1007 900 1009 903
rect 1015 900 1017 903
rect 1105 900 1107 903
rect 1113 900 1115 903
rect 1152 900 1154 903
rect 1160 900 1162 903
rect 1250 900 1252 903
rect 1258 900 1260 903
rect 1297 900 1299 903
rect 1305 900 1307 903
rect 1395 900 1397 903
rect 1403 900 1405 903
rect 1442 900 1444 903
rect 1450 900 1452 903
rect 359 884 368 886
rect 388 884 401 886
rect 421 884 424 886
rect 153 881 165 883
rect 185 881 201 883
rect 221 881 224 883
rect -666 873 -664 876
rect -615 873 -613 876
rect -338 873 -336 876
rect -288 873 -286 876
rect 359 876 368 878
rect 388 876 401 878
rect 421 876 424 878
rect 446 876 448 892
rect 477 883 486 885
rect 526 883 538 885
rect 548 883 551 885
rect 153 873 165 875
rect 185 873 201 875
rect 221 873 224 875
rect 477 875 486 877
rect 526 875 538 877
rect 548 875 551 877
rect 574 876 576 892
rect 446 863 448 866
rect 574 863 576 866
rect 678 864 680 880
rect 686 864 688 880
rect 725 864 727 880
rect 733 864 735 880
rect 820 864 822 880
rect 828 864 830 880
rect 867 864 869 880
rect 875 864 877 880
rect 960 864 962 880
rect 968 864 970 880
rect 1007 864 1009 880
rect 1015 864 1017 880
rect 1105 864 1107 880
rect 1113 864 1115 880
rect 1152 864 1154 880
rect 1160 864 1162 880
rect 1250 864 1252 880
rect 1258 864 1260 880
rect 1297 864 1299 880
rect 1305 864 1307 880
rect 1395 864 1397 880
rect 1403 864 1405 880
rect 1442 864 1444 880
rect 1450 864 1452 880
rect 137 851 139 854
rect 678 832 680 844
rect 686 832 688 844
rect 725 832 727 844
rect 733 832 735 844
rect 820 832 822 844
rect 828 832 830 844
rect 867 832 869 844
rect 875 832 877 844
rect 960 832 962 844
rect 968 832 970 844
rect 1007 832 1009 844
rect 1015 832 1017 844
rect 1105 832 1107 844
rect 1113 832 1115 844
rect 1152 832 1154 844
rect 1160 832 1162 844
rect 1250 832 1252 844
rect 1258 832 1260 844
rect 1297 832 1299 844
rect 1305 832 1307 844
rect 1395 832 1397 844
rect 1403 832 1405 844
rect 1442 832 1444 844
rect 1450 832 1452 844
rect 50 823 59 825
rect 79 823 92 825
rect 112 823 115 825
rect 50 815 59 817
rect 79 815 92 817
rect 112 815 115 817
rect 137 815 139 831
rect 369 826 371 829
rect 522 819 524 822
rect 137 802 139 805
rect 282 798 291 800
rect 311 798 324 800
rect 344 798 347 800
rect 282 790 291 792
rect 311 790 324 792
rect 344 790 347 792
rect 369 790 371 806
rect 406 801 415 803
rect 475 801 487 803
rect 497 801 500 803
rect 702 804 705 806
rect 725 804 739 806
rect 749 804 752 806
rect 844 804 847 806
rect 867 804 881 806
rect 891 804 894 806
rect 984 804 987 806
rect 1007 804 1021 806
rect 1031 804 1034 806
rect 1129 804 1132 806
rect 1152 804 1166 806
rect 1176 804 1179 806
rect 1274 804 1277 806
rect 1297 804 1311 806
rect 1321 804 1324 806
rect 1419 804 1422 806
rect 1442 804 1456 806
rect 1466 804 1469 806
rect 406 793 415 795
rect 475 793 487 795
rect 497 793 500 795
rect 406 785 415 787
rect 475 785 487 787
rect 497 785 500 787
rect 522 783 524 799
rect 369 777 371 780
rect 522 770 524 773
rect 152 757 164 759
rect 184 757 200 759
rect 220 757 223 759
rect 702 753 705 755
rect 725 753 739 755
rect 749 753 752 755
rect 844 753 847 755
rect 867 753 881 755
rect 891 753 894 755
rect 984 753 987 755
rect 1007 753 1021 755
rect 1031 753 1034 755
rect 1129 753 1132 755
rect 1152 753 1166 755
rect 1176 753 1179 755
rect 1274 753 1277 755
rect 1297 753 1311 755
rect 1321 753 1324 755
rect 1419 753 1422 755
rect 1442 753 1456 755
rect 1466 753 1469 755
rect 152 749 164 751
rect 184 749 200 751
rect 220 749 223 751
rect -1140 728 -1128 730
rect -1108 728 -1092 730
rect -1072 728 -1069 730
rect -813 728 -801 730
rect -781 728 -765 730
rect -745 728 -742 730
rect -1140 720 -1128 722
rect -1108 720 -1092 722
rect -1072 720 -1069 722
rect -481 727 -469 729
rect -449 727 -433 729
rect -413 727 -410 729
rect -813 720 -801 722
rect -781 720 -765 722
rect -745 720 -742 722
rect -1246 710 -1234 712
rect -1214 710 -1198 712
rect -1178 710 -1175 712
rect 461 733 463 736
rect -154 727 -142 729
rect -122 727 -106 729
rect -86 727 -83 729
rect -481 719 -469 721
rect -449 719 -433 721
rect -413 719 -410 721
rect -919 710 -907 712
rect -887 710 -871 712
rect -851 710 -848 712
rect -1246 702 -1234 704
rect -1214 702 -1198 704
rect -1178 702 -1175 704
rect 61 723 73 725
rect 93 723 109 725
rect 129 723 132 725
rect -154 719 -142 721
rect -122 719 -106 721
rect -86 719 -83 721
rect -587 709 -575 711
rect -555 709 -539 711
rect -519 709 -516 711
rect -919 702 -907 704
rect -887 702 -871 704
rect -851 702 -848 704
rect 248 723 260 725
rect 280 723 296 725
rect 316 723 319 725
rect 61 715 73 717
rect 93 715 109 717
rect 129 715 132 717
rect -260 709 -248 711
rect -228 709 -212 711
rect -192 709 -189 711
rect 248 715 260 717
rect 280 715 296 717
rect 316 715 319 717
rect 365 716 374 718
rect 394 716 406 718
rect 436 716 439 718
rect -587 701 -575 703
rect -555 701 -539 703
rect -519 701 -516 703
rect -260 701 -248 703
rect -228 701 -212 703
rect -192 701 -189 703
rect 365 708 374 710
rect 394 708 406 710
rect 436 708 439 710
rect 152 701 164 703
rect 184 701 200 703
rect 220 701 223 703
rect 365 700 374 702
rect 394 700 406 702
rect 436 700 439 702
rect 461 697 463 713
rect 152 693 164 695
rect 184 693 200 695
rect 220 693 223 695
rect -1325 685 -1323 688
rect -1274 685 -1272 688
rect -997 685 -995 688
rect -947 685 -945 688
rect -1325 651 -1323 665
rect -1274 651 -1272 665
rect -1246 663 -1234 665
rect -1214 663 -1198 665
rect -1178 663 -1175 665
rect -666 684 -664 687
rect -615 684 -613 687
rect -338 684 -336 687
rect -288 684 -286 687
rect 461 684 463 687
rect -1140 663 -1128 665
rect -1108 663 -1092 665
rect -1072 663 -1069 665
rect -1246 655 -1234 657
rect -1214 655 -1198 657
rect -1178 655 -1175 657
rect -1140 655 -1128 657
rect -1108 655 -1092 657
rect -1072 655 -1069 657
rect -997 651 -995 665
rect -947 651 -945 665
rect -919 663 -907 665
rect -887 663 -871 665
rect -851 663 -848 665
rect -813 663 -801 665
rect -781 663 -765 665
rect -745 663 -742 665
rect -919 655 -907 657
rect -887 655 -871 657
rect -851 655 -848 657
rect -813 655 -801 657
rect -781 655 -765 657
rect -745 655 -742 657
rect -666 650 -664 664
rect -615 650 -613 664
rect -587 662 -575 664
rect -555 662 -539 664
rect -519 662 -516 664
rect 136 671 138 674
rect -481 662 -469 664
rect -449 662 -433 664
rect -413 662 -410 664
rect -587 654 -575 656
rect -555 654 -539 656
rect -519 654 -516 656
rect -1325 638 -1323 641
rect -1274 638 -1272 641
rect -997 638 -995 641
rect -947 638 -945 641
rect -481 654 -469 656
rect -449 654 -433 656
rect -413 654 -410 656
rect -338 650 -336 664
rect -288 650 -286 664
rect -260 662 -248 664
rect -228 662 -212 664
rect -192 662 -189 664
rect -154 662 -142 664
rect -122 662 -106 664
rect -86 662 -83 664
rect -260 654 -248 656
rect -228 654 -212 656
rect -192 654 -189 656
rect -154 654 -142 656
rect -122 654 -106 656
rect -86 654 -83 656
rect 643 670 655 672
rect 675 670 691 672
rect 711 670 714 672
rect 643 662 655 664
rect 675 662 691 664
rect 711 662 714 664
rect 49 643 58 645
rect 78 643 91 645
rect 111 643 114 645
rect -666 637 -664 640
rect -615 637 -613 640
rect -338 637 -336 640
rect -288 637 -286 640
rect 49 635 58 637
rect 78 635 91 637
rect 111 635 114 637
rect 136 635 138 651
rect 552 636 564 638
rect 584 636 600 638
rect 620 636 623 638
rect 284 630 296 632
rect 316 630 332 632
rect 352 630 355 632
rect 136 622 138 625
rect 739 636 751 638
rect 771 636 787 638
rect 807 636 810 638
rect 552 628 564 630
rect 584 628 600 630
rect 620 628 623 630
rect 284 622 296 624
rect 316 622 332 624
rect 352 622 355 624
rect 739 628 751 630
rect 771 628 787 630
rect 807 628 810 630
rect 643 614 655 616
rect 675 614 691 616
rect 711 614 714 616
rect 643 606 655 608
rect 675 606 691 608
rect 711 606 714 608
rect 193 596 205 598
rect 225 596 241 598
rect 261 596 264 598
rect 380 596 392 598
rect 412 596 428 598
rect 448 596 451 598
rect 193 588 205 590
rect 225 588 241 590
rect 261 588 264 590
rect 380 588 392 590
rect 412 588 428 590
rect 448 588 451 590
rect 284 574 296 576
rect 316 574 332 576
rect 352 574 355 576
rect 284 566 296 568
rect 316 566 332 568
rect 352 566 355 568
rect 626 560 628 563
rect 539 532 548 534
rect 568 532 581 534
rect 601 532 604 534
rect 539 524 548 526
rect 568 524 581 526
rect 601 524 604 526
rect 626 524 628 540
rect -1140 514 -1128 516
rect -1108 514 -1092 516
rect -1072 514 -1069 516
rect -813 514 -801 516
rect -781 514 -765 516
rect -745 514 -742 516
rect -1140 506 -1128 508
rect -1108 506 -1092 508
rect -1072 506 -1069 508
rect -481 513 -469 515
rect -449 513 -433 515
rect -413 513 -410 515
rect -813 506 -801 508
rect -781 506 -765 508
rect -745 506 -742 508
rect -1246 496 -1234 498
rect -1214 496 -1198 498
rect -1178 496 -1175 498
rect -154 513 -142 515
rect -122 513 -106 515
rect -86 513 -83 515
rect -481 505 -469 507
rect -449 505 -433 507
rect -413 505 -410 507
rect -919 496 -907 498
rect -887 496 -871 498
rect -851 496 -848 498
rect -1246 488 -1234 490
rect -1214 488 -1198 490
rect -1178 488 -1175 490
rect 626 511 628 514
rect -154 505 -142 507
rect -122 505 -106 507
rect -86 505 -83 507
rect -587 495 -575 497
rect -555 495 -539 497
rect -519 495 -516 497
rect -919 488 -907 490
rect -887 488 -871 490
rect -851 488 -848 490
rect 823 507 825 510
rect 152 503 164 505
rect 184 503 200 505
rect 220 503 223 505
rect -260 495 -248 497
rect -228 495 -212 497
rect -192 495 -189 497
rect -587 487 -575 489
rect -555 487 -539 489
rect -519 487 -516 489
rect 152 495 164 497
rect 184 495 200 497
rect 220 495 223 497
rect 476 495 478 498
rect 635 496 637 499
rect -260 487 -248 489
rect -228 487 -212 489
rect -192 487 -189 489
rect 370 481 379 483
rect 399 481 411 483
rect 451 481 454 483
rect -1325 471 -1323 474
rect -1274 471 -1272 474
rect -997 471 -995 474
rect -947 471 -945 474
rect -1325 437 -1323 451
rect -1274 437 -1272 451
rect -1246 449 -1234 451
rect -1214 449 -1198 451
rect -1178 449 -1175 451
rect -666 470 -664 473
rect -615 470 -613 473
rect -338 470 -336 473
rect -288 470 -286 473
rect -1140 449 -1128 451
rect -1108 449 -1092 451
rect -1072 449 -1069 451
rect -1246 441 -1234 443
rect -1214 441 -1198 443
rect -1178 441 -1175 443
rect -1140 441 -1128 443
rect -1108 441 -1092 443
rect -1072 441 -1069 443
rect -997 437 -995 451
rect -947 437 -945 451
rect -919 449 -907 451
rect -887 449 -871 451
rect -851 449 -848 451
rect -813 449 -801 451
rect -781 449 -765 451
rect -745 449 -742 451
rect -919 441 -907 443
rect -887 441 -871 443
rect -851 441 -848 443
rect -813 441 -801 443
rect -781 441 -765 443
rect -745 441 -742 443
rect -666 436 -664 450
rect -615 436 -613 450
rect -587 448 -575 450
rect -555 448 -539 450
rect -519 448 -516 450
rect 61 469 73 471
rect 93 469 109 471
rect 129 469 132 471
rect 539 479 548 481
rect 568 479 580 481
rect 610 479 613 481
rect 370 473 379 475
rect 399 473 411 475
rect 451 473 454 475
rect 248 469 260 471
rect 280 469 296 471
rect 316 469 319 471
rect 61 461 73 463
rect 93 461 109 463
rect 129 461 132 463
rect 370 465 379 467
rect 399 465 411 467
rect 451 465 454 467
rect 248 461 260 463
rect 280 461 296 463
rect 316 461 319 463
rect 476 459 478 475
rect 686 495 695 497
rect 775 495 787 497
rect 797 495 800 497
rect 686 487 695 489
rect 775 487 787 489
rect 797 487 800 489
rect 686 479 695 481
rect 775 479 787 481
rect 797 479 800 481
rect 539 471 548 473
rect 568 471 580 473
rect 610 471 613 473
rect 539 463 548 465
rect 568 463 580 465
rect 610 463 613 465
rect 370 457 379 459
rect 399 457 411 459
rect 451 457 454 459
rect -481 448 -469 450
rect -449 448 -433 450
rect -413 448 -410 450
rect -587 440 -575 442
rect -555 440 -539 442
rect -519 440 -516 442
rect -1325 424 -1323 427
rect -1274 424 -1272 427
rect -997 424 -995 427
rect -947 424 -945 427
rect -481 440 -469 442
rect -449 440 -433 442
rect -413 440 -410 442
rect -338 436 -336 450
rect -288 436 -286 450
rect -260 448 -248 450
rect -228 448 -212 450
rect -192 448 -189 450
rect -154 448 -142 450
rect -122 448 -106 450
rect -86 448 -83 450
rect -260 440 -248 442
rect -228 440 -212 442
rect -192 440 -189 442
rect 635 460 637 476
rect 686 471 695 473
rect 775 471 787 473
rect 797 471 800 473
rect 823 471 825 487
rect 823 458 825 461
rect 152 447 164 449
rect 184 447 200 449
rect 220 447 223 449
rect -154 440 -142 442
rect -122 440 -106 442
rect -86 440 -83 442
rect 476 446 478 449
rect 635 447 637 450
rect 152 439 164 441
rect 184 439 200 441
rect 220 439 223 441
rect 803 439 805 442
rect -666 423 -664 426
rect -615 423 -613 426
rect -338 423 -336 426
rect -288 423 -286 426
rect 136 417 138 420
rect 716 411 725 413
rect 745 411 758 413
rect 778 411 781 413
rect 716 403 725 405
rect 745 403 758 405
rect 778 403 781 405
rect 803 403 805 419
rect 49 389 58 391
rect 78 389 91 391
rect 111 389 114 391
rect 49 381 58 383
rect 78 381 91 383
rect 111 381 114 383
rect 136 381 138 397
rect 803 390 805 393
rect 390 383 392 386
rect 540 384 542 387
rect 676 384 678 387
rect 136 368 138 371
rect 298 368 307 370
rect 327 368 339 370
rect 364 368 367 370
rect 434 370 443 372
rect 463 370 475 372
rect 515 370 518 372
rect 298 360 307 362
rect 327 360 339 362
rect 364 360 367 362
rect 298 352 307 354
rect 327 352 339 354
rect 364 352 367 354
rect 390 347 392 363
rect 580 367 589 369
rect 609 367 621 369
rect 651 367 654 369
rect 434 362 443 364
rect 463 362 475 364
rect 515 362 518 364
rect 434 354 443 356
rect 463 354 475 356
rect 515 354 518 356
rect 298 344 307 346
rect 327 344 339 346
rect 364 344 377 346
rect 375 341 377 344
rect 298 336 307 338
rect 327 336 339 338
rect 364 336 367 338
rect 540 348 542 364
rect 580 359 589 361
rect 609 359 621 361
rect 651 359 654 361
rect 580 351 589 353
rect 609 351 621 353
rect 651 351 654 353
rect 434 346 443 348
rect 463 346 475 348
rect 515 346 518 348
rect 676 348 678 364
rect 881 363 883 366
rect 726 347 735 349
rect 835 347 847 349
rect 857 347 860 349
rect 726 339 735 341
rect 835 339 847 341
rect 857 339 860 341
rect 390 334 392 337
rect 540 335 542 338
rect 676 335 678 338
rect 726 331 735 333
rect 835 331 847 333
rect 857 331 860 333
rect 153 321 165 323
rect 185 321 201 323
rect 221 321 224 323
rect 881 327 883 343
rect 726 323 735 325
rect 835 323 847 325
rect 857 323 860 325
rect 153 313 165 315
rect 185 313 201 315
rect 221 313 224 315
rect 726 315 735 317
rect 835 315 847 317
rect 857 315 860 317
rect 881 314 883 317
rect 62 287 74 289
rect 94 287 110 289
rect 130 287 133 289
rect -1140 275 -1128 277
rect -1108 275 -1092 277
rect -1072 275 -1069 277
rect -813 275 -801 277
rect -781 275 -765 277
rect -745 275 -742 277
rect -1140 267 -1128 269
rect -1108 267 -1092 269
rect -1072 267 -1069 269
rect -481 274 -469 276
rect -449 274 -433 276
rect -413 274 -410 276
rect -813 267 -801 269
rect -781 267 -765 269
rect -745 267 -742 269
rect -1246 257 -1234 259
rect -1214 257 -1198 259
rect -1178 257 -1175 259
rect 249 287 261 289
rect 281 287 297 289
rect 317 287 320 289
rect 62 279 74 281
rect 94 279 110 281
rect 130 279 133 281
rect -154 274 -142 276
rect -122 274 -106 276
rect -86 274 -83 276
rect 249 279 261 281
rect 281 279 297 281
rect 317 279 320 281
rect -481 266 -469 268
rect -449 266 -433 268
rect -413 266 -410 268
rect -919 257 -907 259
rect -887 257 -871 259
rect -851 257 -848 259
rect -1246 249 -1234 251
rect -1214 249 -1198 251
rect -1178 249 -1175 251
rect -154 266 -142 268
rect -122 266 -106 268
rect -86 266 -83 268
rect -587 256 -575 258
rect -555 256 -539 258
rect -519 256 -516 258
rect -919 249 -907 251
rect -887 249 -871 251
rect -851 249 -848 251
rect 153 265 165 267
rect 185 265 201 267
rect 221 265 224 267
rect -260 256 -248 258
rect -228 256 -212 258
rect -192 256 -189 258
rect 153 257 165 259
rect 185 257 201 259
rect 221 257 224 259
rect -587 248 -575 250
rect -555 248 -539 250
rect -519 248 -516 250
rect 476 252 488 254
rect 508 252 524 254
rect 544 252 547 254
rect -260 248 -248 250
rect -228 248 -212 250
rect -192 248 -189 250
rect 1101 249 1113 251
rect 1133 249 1149 251
rect 1169 249 1172 251
rect 476 244 488 246
rect 508 244 524 246
rect 544 244 547 246
rect 930 239 932 242
rect 1101 241 1113 243
rect 1133 241 1149 243
rect 1169 241 1172 243
rect 137 235 139 238
rect -1325 232 -1323 235
rect -1274 232 -1272 235
rect -997 232 -995 235
rect -947 232 -945 235
rect -1325 198 -1323 212
rect -1274 198 -1272 212
rect -1246 210 -1234 212
rect -1214 210 -1198 212
rect -1178 210 -1175 212
rect -666 231 -664 234
rect -615 231 -613 234
rect -338 231 -336 234
rect -288 231 -286 234
rect -1140 210 -1128 212
rect -1108 210 -1092 212
rect -1072 210 -1069 212
rect -1246 202 -1234 204
rect -1214 202 -1198 204
rect -1178 202 -1175 204
rect -1140 202 -1128 204
rect -1108 202 -1092 204
rect -1072 202 -1069 204
rect -997 198 -995 212
rect -947 198 -945 212
rect -919 210 -907 212
rect -887 210 -871 212
rect -851 210 -848 212
rect -813 210 -801 212
rect -781 210 -765 212
rect -745 210 -742 212
rect -919 202 -907 204
rect -887 202 -871 204
rect -851 202 -848 204
rect -813 202 -801 204
rect -781 202 -765 204
rect -745 202 -742 204
rect -666 197 -664 211
rect -615 197 -613 211
rect -587 209 -575 211
rect -555 209 -539 211
rect -519 209 -516 211
rect -481 209 -469 211
rect -449 209 -433 211
rect -413 209 -410 211
rect -587 201 -575 203
rect -555 201 -539 203
rect -519 201 -516 203
rect -1325 185 -1323 188
rect -1274 185 -1272 188
rect -997 185 -995 188
rect -947 185 -945 188
rect -481 201 -469 203
rect -449 201 -433 203
rect -413 201 -410 203
rect -338 197 -336 211
rect -288 197 -286 211
rect -260 209 -248 211
rect -228 209 -212 211
rect -192 209 -189 211
rect 385 218 397 220
rect 417 218 433 220
rect 453 218 456 220
rect -154 209 -142 211
rect -122 209 -106 211
rect -86 209 -83 211
rect -260 201 -248 203
rect -228 201 -212 203
rect -192 201 -189 203
rect 50 207 59 209
rect 79 207 92 209
rect 112 207 115 209
rect -154 201 -142 203
rect -122 201 -106 203
rect -86 201 -83 203
rect 50 199 59 201
rect 79 199 92 201
rect 112 199 115 201
rect 137 199 139 215
rect 572 218 584 220
rect 604 218 620 220
rect 640 218 643 220
rect 385 210 397 212
rect 417 210 433 212
rect 453 210 456 212
rect 793 216 795 219
rect 572 210 584 212
rect 604 210 620 212
rect 640 210 643 212
rect 697 199 706 201
rect 726 199 738 201
rect 768 199 771 201
rect 476 196 488 198
rect 508 196 524 198
rect 544 196 547 198
rect -666 184 -664 187
rect -615 184 -613 187
rect -338 184 -336 187
rect -288 184 -286 187
rect 137 186 139 189
rect 843 211 852 213
rect 872 211 885 213
rect 905 211 908 213
rect 843 203 852 205
rect 872 203 885 205
rect 905 203 908 205
rect 930 203 932 219
rect 1010 215 1022 217
rect 1042 215 1058 217
rect 1078 215 1081 217
rect 1197 215 1209 217
rect 1229 215 1245 217
rect 1265 215 1268 217
rect 1010 207 1022 209
rect 1042 207 1058 209
rect 1078 207 1081 209
rect 697 191 706 193
rect 726 191 738 193
rect 768 191 771 193
rect 476 188 488 190
rect 508 188 524 190
rect 544 188 547 190
rect 697 183 706 185
rect 726 183 738 185
rect 768 183 771 185
rect 793 180 795 196
rect 1197 207 1209 209
rect 1229 207 1245 209
rect 1265 207 1268 209
rect 930 190 932 193
rect 1101 193 1113 195
rect 1133 193 1149 195
rect 1169 193 1172 195
rect 1101 185 1113 187
rect 1133 185 1149 187
rect 1169 185 1172 187
rect 793 167 795 170
rect 608 145 610 148
rect 154 138 166 140
rect 186 138 202 140
rect 222 138 225 140
rect 475 136 477 139
rect 154 130 166 132
rect 186 130 202 132
rect 222 130 225 132
rect 379 128 389 130
rect 399 128 413 130
rect 443 128 446 130
rect 379 120 389 122
rect 399 120 413 122
rect 443 120 446 122
rect 516 130 525 132
rect 545 130 557 132
rect 582 130 585 132
rect 750 136 752 139
rect 516 122 525 124
rect 545 122 557 124
rect 582 122 585 124
rect 379 112 389 114
rect 399 112 413 114
rect 443 112 446 114
rect 63 104 75 106
rect 95 104 111 106
rect 131 104 134 106
rect 250 104 262 106
rect 282 104 298 106
rect 318 104 321 106
rect 63 96 75 98
rect 95 96 111 98
rect 131 96 134 98
rect -1140 88 -1128 90
rect -1108 88 -1092 90
rect -1072 88 -1069 90
rect -813 88 -801 90
rect -781 88 -765 90
rect -745 88 -742 90
rect -1140 80 -1128 82
rect -1108 80 -1092 82
rect -1072 80 -1069 82
rect -481 87 -469 89
rect -449 87 -433 89
rect -413 87 -410 89
rect -813 80 -801 82
rect -781 80 -765 82
rect -745 80 -742 82
rect -1246 70 -1234 72
rect -1214 70 -1198 72
rect -1178 70 -1175 72
rect 379 104 389 106
rect 399 104 413 106
rect 443 104 446 106
rect 250 96 262 98
rect 282 96 298 98
rect 318 96 321 98
rect 475 100 477 116
rect 516 114 525 116
rect 545 114 557 116
rect 582 114 585 116
rect 608 109 610 125
rect 644 122 653 124
rect 673 122 685 124
rect 725 122 728 124
rect 1039 134 1041 137
rect 853 126 864 128
rect 984 126 996 128
rect 1006 126 1009 128
rect 853 118 864 120
rect 984 118 996 120
rect 1006 118 1009 120
rect 644 114 653 116
rect 673 114 685 116
rect 725 114 728 116
rect 516 106 525 108
rect 545 106 557 108
rect 582 106 597 108
rect 379 96 389 98
rect 399 96 413 98
rect 443 96 446 98
rect -154 87 -142 89
rect -122 87 -106 89
rect -86 87 -83 89
rect -481 79 -469 81
rect -449 79 -433 81
rect -413 79 -410 81
rect -919 70 -907 72
rect -887 70 -871 72
rect -851 70 -848 72
rect -1246 62 -1234 64
rect -1214 62 -1198 64
rect -1178 62 -1175 64
rect 516 98 525 100
rect 545 98 557 100
rect 582 98 585 100
rect 644 106 653 108
rect 673 106 685 108
rect 725 106 728 108
rect 608 96 610 99
rect 750 100 752 116
rect 853 110 864 112
rect 984 110 996 112
rect 1006 110 1009 112
rect 853 102 864 104
rect 984 102 996 104
rect 1006 102 1009 104
rect 644 98 653 100
rect 673 98 685 100
rect 725 98 728 100
rect 1039 98 1041 114
rect 853 94 864 96
rect 984 94 996 96
rect 1006 94 1009 96
rect 379 88 389 90
rect 399 88 413 90
rect 443 88 446 90
rect 154 82 166 84
rect 186 82 202 84
rect 222 82 225 84
rect 475 87 477 90
rect 750 87 752 90
rect 853 86 864 88
rect 984 86 996 88
rect 1006 86 1009 88
rect -154 79 -142 81
rect -122 79 -106 81
rect -86 79 -83 81
rect -587 69 -575 71
rect -555 69 -539 71
rect -519 69 -516 71
rect -919 62 -907 64
rect -887 62 -871 64
rect -851 62 -848 64
rect 1039 85 1041 88
rect 154 74 166 76
rect 186 74 202 76
rect 222 74 225 76
rect -260 69 -248 71
rect -228 69 -212 71
rect -192 69 -189 71
rect -587 61 -575 63
rect -555 61 -539 63
rect -519 61 -516 63
rect -260 61 -248 63
rect -228 61 -212 63
rect -192 61 -189 63
rect 138 52 140 55
rect -1325 45 -1323 48
rect -1274 45 -1272 48
rect -997 45 -995 48
rect -947 45 -945 48
rect -1325 11 -1323 25
rect -1274 11 -1272 25
rect -1246 23 -1234 25
rect -1214 23 -1198 25
rect -1178 23 -1175 25
rect -666 44 -664 47
rect -615 44 -613 47
rect -338 44 -336 47
rect -288 44 -286 47
rect -1140 23 -1128 25
rect -1108 23 -1092 25
rect -1072 23 -1069 25
rect -1246 15 -1234 17
rect -1214 15 -1198 17
rect -1178 15 -1175 17
rect -1140 15 -1128 17
rect -1108 15 -1092 17
rect -1072 15 -1069 17
rect -997 11 -995 25
rect -947 11 -945 25
rect -919 23 -907 25
rect -887 23 -871 25
rect -851 23 -848 25
rect -813 23 -801 25
rect -781 23 -765 25
rect -745 23 -742 25
rect -919 15 -907 17
rect -887 15 -871 17
rect -851 15 -848 17
rect -813 15 -801 17
rect -781 15 -765 17
rect -745 15 -742 17
rect -666 10 -664 24
rect -615 10 -613 24
rect -587 22 -575 24
rect -555 22 -539 24
rect -519 22 -516 24
rect -481 22 -469 24
rect -449 22 -433 24
rect -413 22 -410 24
rect -587 14 -575 16
rect -555 14 -539 16
rect -519 14 -516 16
rect -1325 -2 -1323 1
rect -1274 -2 -1272 1
rect -997 -2 -995 1
rect -947 -2 -945 1
rect -481 14 -469 16
rect -449 14 -433 16
rect -413 14 -410 16
rect -338 10 -336 24
rect -288 10 -286 24
rect -260 22 -248 24
rect -228 22 -212 24
rect -192 22 -189 24
rect -154 22 -142 24
rect -122 22 -106 24
rect -86 22 -83 24
rect 51 24 60 26
rect 80 24 93 26
rect 113 24 116 26
rect -260 14 -248 16
rect -228 14 -212 16
rect -192 14 -189 16
rect -154 14 -142 16
rect -122 14 -106 16
rect -86 14 -83 16
rect 51 16 60 18
rect 80 16 93 18
rect 113 16 116 18
rect 138 16 140 32
rect 138 3 140 6
rect -666 -3 -664 0
rect -615 -3 -613 0
rect -338 -3 -336 0
rect -288 -3 -286 0
<< ndiffusion >>
rect 659 1313 660 1333
rect 662 1313 663 1333
rect 667 1313 668 1333
rect 670 1313 671 1333
rect 724 1313 725 1333
rect 727 1313 728 1333
rect 732 1313 733 1333
rect 735 1313 736 1333
rect 801 1313 802 1333
rect 804 1313 805 1333
rect 809 1313 810 1333
rect 812 1313 813 1333
rect 866 1313 867 1333
rect 869 1313 870 1333
rect 874 1313 875 1333
rect 877 1313 878 1333
rect 941 1313 942 1333
rect 944 1313 945 1333
rect 949 1313 950 1333
rect 952 1313 953 1333
rect 1006 1313 1007 1333
rect 1009 1313 1010 1333
rect 1014 1313 1015 1333
rect 1017 1313 1018 1333
rect 1086 1313 1087 1333
rect 1089 1313 1090 1333
rect 1094 1313 1095 1333
rect 1097 1313 1098 1333
rect 1151 1313 1152 1333
rect 1154 1313 1155 1333
rect 1159 1313 1160 1333
rect 1162 1313 1163 1333
rect 1231 1313 1232 1333
rect 1234 1313 1235 1333
rect 1239 1313 1240 1333
rect 1242 1313 1243 1333
rect 1296 1313 1297 1333
rect 1299 1313 1300 1333
rect 1304 1313 1305 1333
rect 1307 1313 1308 1333
rect 1376 1313 1377 1333
rect 1379 1313 1380 1333
rect 1384 1313 1385 1333
rect 1387 1313 1388 1333
rect 1441 1313 1442 1333
rect 1444 1313 1445 1333
rect 1449 1313 1450 1333
rect 1452 1313 1453 1333
rect 677 1207 678 1227
rect 680 1207 681 1227
rect 685 1207 686 1227
rect 688 1207 689 1227
rect 724 1207 725 1227
rect 727 1207 728 1227
rect 732 1207 733 1227
rect 735 1207 736 1227
rect 819 1207 820 1227
rect 822 1207 823 1227
rect 827 1207 828 1227
rect 830 1207 831 1227
rect 866 1207 867 1227
rect 869 1207 870 1227
rect 874 1207 875 1227
rect 877 1207 878 1227
rect 959 1207 960 1227
rect 962 1207 963 1227
rect 967 1207 968 1227
rect 970 1207 971 1227
rect 1006 1207 1007 1227
rect 1009 1207 1010 1227
rect 1014 1207 1015 1227
rect 1017 1207 1018 1227
rect 1104 1207 1105 1227
rect 1107 1207 1108 1227
rect 1112 1207 1113 1227
rect 1115 1207 1116 1227
rect 1151 1207 1152 1227
rect 1154 1207 1155 1227
rect 1159 1207 1160 1227
rect 1162 1207 1163 1227
rect 1249 1207 1250 1227
rect 1252 1207 1253 1227
rect 1257 1207 1258 1227
rect 1260 1207 1261 1227
rect 1296 1207 1297 1227
rect 1299 1207 1300 1227
rect 1304 1207 1305 1227
rect 1307 1207 1308 1227
rect 1394 1207 1395 1227
rect 1397 1207 1398 1227
rect 1402 1207 1403 1227
rect 1405 1207 1406 1227
rect 1441 1207 1442 1227
rect 1444 1207 1445 1227
rect 1449 1207 1450 1227
rect 1452 1207 1453 1227
rect -432 1129 -412 1130
rect -432 1126 -412 1127
rect 739 1133 749 1134
rect 881 1133 891 1134
rect 1021 1133 1031 1134
rect 1166 1133 1176 1134
rect 1311 1133 1321 1134
rect 1456 1133 1466 1134
rect -105 1129 -85 1130
rect -432 1121 -412 1122
rect -432 1118 -412 1119
rect -105 1126 -85 1127
rect 739 1130 749 1131
rect 881 1130 891 1131
rect 1021 1130 1031 1131
rect 1166 1130 1176 1131
rect 1311 1130 1321 1131
rect 1456 1130 1466 1131
rect -105 1121 -85 1122
rect -538 1111 -518 1112
rect -538 1108 -518 1109
rect -105 1118 -85 1119
rect -211 1111 -191 1112
rect -538 1103 -518 1104
rect -538 1100 -518 1101
rect -211 1108 -191 1109
rect -211 1103 -191 1104
rect -211 1100 -191 1101
rect -538 1064 -518 1065
rect -538 1061 -518 1062
rect -432 1064 -412 1065
rect 739 1083 749 1084
rect 881 1083 891 1084
rect 1021 1083 1031 1084
rect 1166 1083 1176 1084
rect 1311 1083 1321 1084
rect 1456 1083 1466 1084
rect 739 1080 749 1081
rect 881 1080 891 1081
rect 1021 1080 1031 1081
rect 1166 1080 1176 1081
rect 1311 1080 1321 1081
rect 1456 1080 1466 1081
rect -538 1056 -518 1057
rect -666 1040 -665 1050
rect -663 1040 -662 1050
rect -615 1040 -614 1050
rect -612 1040 -611 1050
rect -538 1053 -518 1054
rect -432 1061 -412 1062
rect -432 1056 -412 1057
rect -432 1053 -412 1054
rect -211 1064 -191 1065
rect -211 1061 -191 1062
rect -105 1064 -85 1065
rect -211 1056 -191 1057
rect -338 1040 -337 1050
rect -335 1040 -334 1050
rect -288 1040 -287 1050
rect -285 1040 -284 1050
rect -211 1053 -191 1054
rect -105 1061 -85 1062
rect -105 1056 -85 1057
rect -105 1053 -85 1054
rect 452 1027 472 1028
rect 452 1024 472 1025
rect 452 1019 472 1020
rect 452 1016 472 1017
rect 361 993 381 994
rect 361 990 381 991
rect 548 993 568 994
rect 361 985 381 986
rect 361 982 381 983
rect 548 990 568 991
rect 659 986 660 1006
rect 662 986 663 1006
rect 667 986 668 1006
rect 670 986 671 1006
rect 724 986 725 1006
rect 727 986 728 1006
rect 732 986 733 1006
rect 735 986 736 1006
rect 801 986 802 1006
rect 804 986 805 1006
rect 809 986 810 1006
rect 812 986 813 1006
rect 866 986 867 1006
rect 869 986 870 1006
rect 874 986 875 1006
rect 877 986 878 1006
rect 941 986 942 1006
rect 944 986 945 1006
rect 949 986 950 1006
rect 952 986 953 1006
rect 1006 986 1007 1006
rect 1009 986 1010 1006
rect 1014 986 1015 1006
rect 1017 986 1018 1006
rect 1086 986 1087 1006
rect 1089 986 1090 1006
rect 1094 986 1095 1006
rect 1097 986 1098 1006
rect 1151 986 1152 1006
rect 1154 986 1155 1006
rect 1159 986 1160 1006
rect 1162 986 1163 1006
rect 1231 986 1232 1006
rect 1234 986 1235 1006
rect 1239 986 1240 1006
rect 1242 986 1243 1006
rect 1296 986 1297 1006
rect 1299 986 1300 1006
rect 1304 986 1305 1006
rect 1307 986 1308 1006
rect 1376 986 1377 1006
rect 1379 986 1380 1006
rect 1384 986 1385 1006
rect 1387 986 1388 1006
rect 1441 986 1442 1006
rect 1444 986 1445 1006
rect 1449 986 1450 1006
rect 1452 986 1453 1006
rect 548 985 568 986
rect 548 982 568 983
rect -1092 969 -1072 970
rect -1092 966 -1072 967
rect -765 969 -745 970
rect -1092 961 -1072 962
rect -1092 958 -1072 959
rect -765 966 -745 967
rect -433 965 -413 966
rect -765 961 -745 962
rect -1198 951 -1178 952
rect -1198 948 -1178 949
rect -765 958 -745 959
rect -433 962 -413 963
rect 452 971 472 972
rect -106 965 -86 966
rect -433 957 -413 958
rect -871 951 -851 952
rect -1198 943 -1178 944
rect -1198 940 -1178 941
rect -871 948 -851 949
rect -433 954 -413 955
rect -106 962 -86 963
rect 452 968 472 969
rect 452 963 472 964
rect -106 957 -86 958
rect 452 960 472 961
rect -539 947 -519 948
rect -871 943 -851 944
rect -871 940 -851 941
rect -539 944 -519 945
rect -106 954 -86 955
rect -212 947 -192 948
rect -539 939 -519 940
rect -539 936 -519 937
rect -212 944 -192 945
rect -212 939 -192 940
rect -212 936 -192 937
rect 201 939 221 940
rect 201 936 221 937
rect 201 931 221 932
rect 201 928 221 929
rect -1198 904 -1178 905
rect -1198 901 -1178 902
rect -1092 904 -1072 905
rect -1198 896 -1178 897
rect -1326 880 -1325 890
rect -1323 880 -1322 890
rect -1275 880 -1274 890
rect -1272 880 -1271 890
rect -1198 893 -1178 894
rect -1092 901 -1072 902
rect -1092 896 -1072 897
rect -1092 893 -1072 894
rect -871 904 -851 905
rect -871 901 -851 902
rect -765 904 -745 905
rect -871 896 -851 897
rect -998 880 -997 890
rect -995 880 -994 890
rect -948 880 -947 890
rect -945 880 -944 890
rect -871 893 -851 894
rect -765 901 -745 902
rect -765 896 -745 897
rect -765 893 -745 894
rect -539 900 -519 901
rect -539 897 -519 898
rect -433 900 -413 901
rect -539 892 -519 893
rect -667 876 -666 886
rect -664 876 -663 886
rect -616 876 -615 886
rect -613 876 -612 886
rect -539 889 -519 890
rect -433 897 -413 898
rect -433 892 -413 893
rect -433 889 -413 890
rect -212 900 -192 901
rect -212 897 -192 898
rect 110 905 130 906
rect -106 900 -86 901
rect -212 892 -192 893
rect -339 876 -338 886
rect -336 876 -335 886
rect -289 876 -288 886
rect -286 876 -285 886
rect -212 889 -192 890
rect -106 897 -86 898
rect 110 902 130 903
rect 297 905 317 906
rect 110 897 130 898
rect -106 892 -86 893
rect 110 894 130 895
rect 297 902 317 903
rect 297 897 317 898
rect 297 894 317 895
rect -106 889 -86 890
rect 201 883 221 884
rect 401 886 421 887
rect 201 880 221 881
rect 201 875 221 876
rect 401 883 421 884
rect 401 878 421 879
rect 538 885 548 886
rect 201 872 221 873
rect 401 875 421 876
rect 445 866 446 876
rect 448 866 449 876
rect 538 882 548 883
rect 538 877 548 878
rect 677 880 678 900
rect 680 880 681 900
rect 685 880 686 900
rect 688 880 689 900
rect 724 880 725 900
rect 727 880 728 900
rect 732 880 733 900
rect 735 880 736 900
rect 819 880 820 900
rect 822 880 823 900
rect 827 880 828 900
rect 830 880 831 900
rect 866 880 867 900
rect 869 880 870 900
rect 874 880 875 900
rect 877 880 878 900
rect 959 880 960 900
rect 962 880 963 900
rect 967 880 968 900
rect 970 880 971 900
rect 1006 880 1007 900
rect 1009 880 1010 900
rect 1014 880 1015 900
rect 1017 880 1018 900
rect 1104 880 1105 900
rect 1107 880 1108 900
rect 1112 880 1113 900
rect 1115 880 1116 900
rect 1151 880 1152 900
rect 1154 880 1155 900
rect 1159 880 1160 900
rect 1162 880 1163 900
rect 1249 880 1250 900
rect 1252 880 1253 900
rect 1257 880 1258 900
rect 1260 880 1261 900
rect 1296 880 1297 900
rect 1299 880 1300 900
rect 1304 880 1305 900
rect 1307 880 1308 900
rect 1394 880 1395 900
rect 1397 880 1398 900
rect 1402 880 1403 900
rect 1405 880 1406 900
rect 1441 880 1442 900
rect 1444 880 1445 900
rect 1449 880 1450 900
rect 1452 880 1453 900
rect 538 874 548 875
rect 573 866 574 876
rect 576 866 577 876
rect 92 825 112 826
rect 92 822 112 823
rect 92 817 112 818
rect 92 814 112 815
rect 136 805 137 815
rect 139 805 140 815
rect 324 800 344 801
rect 324 797 344 798
rect 324 792 344 793
rect 487 803 497 804
rect 487 800 497 801
rect 739 806 749 807
rect 881 806 891 807
rect 1021 806 1031 807
rect 1166 806 1176 807
rect 1311 806 1321 807
rect 1456 806 1466 807
rect 739 803 749 804
rect 881 803 891 804
rect 1021 803 1031 804
rect 1166 803 1176 804
rect 1311 803 1321 804
rect 1456 803 1466 804
rect 487 795 497 796
rect 324 789 344 790
rect 368 780 369 790
rect 371 780 372 790
rect 487 792 497 793
rect 487 787 497 788
rect 487 784 497 785
rect 521 773 522 783
rect 524 773 525 783
rect 200 759 220 760
rect 200 756 220 757
rect 739 755 749 756
rect 881 755 891 756
rect 1021 755 1031 756
rect 1166 755 1176 756
rect 1311 755 1321 756
rect 1456 755 1466 756
rect 200 751 220 752
rect 200 748 220 749
rect 739 752 749 753
rect 881 752 891 753
rect 1021 752 1031 753
rect 1166 752 1176 753
rect 1311 752 1321 753
rect 1456 752 1466 753
rect -1092 730 -1072 731
rect -1092 727 -1072 728
rect -765 730 -745 731
rect -1092 722 -1072 723
rect -1092 719 -1072 720
rect -765 727 -745 728
rect -433 729 -413 730
rect -765 722 -745 723
rect -1198 712 -1178 713
rect -1198 709 -1178 710
rect -765 719 -745 720
rect -433 726 -413 727
rect -106 729 -86 730
rect -433 721 -413 722
rect -871 712 -851 713
rect -1198 704 -1178 705
rect -1198 701 -1178 702
rect -871 709 -851 710
rect -433 718 -413 719
rect -106 726 -86 727
rect 109 725 129 726
rect -106 721 -86 722
rect -539 711 -519 712
rect -871 704 -851 705
rect -871 701 -851 702
rect -539 708 -519 709
rect -106 718 -86 719
rect 109 722 129 723
rect 296 725 316 726
rect 109 717 129 718
rect -212 711 -192 712
rect 109 714 129 715
rect 296 722 316 723
rect 296 717 316 718
rect 406 718 436 719
rect 296 714 316 715
rect -539 703 -519 704
rect -539 700 -519 701
rect -212 708 -192 709
rect -212 703 -192 704
rect -212 700 -192 701
rect 406 715 436 716
rect 406 710 436 711
rect 200 703 220 704
rect 200 700 220 701
rect 406 707 436 708
rect 406 702 436 703
rect 200 695 220 696
rect 406 699 436 700
rect 200 692 220 693
rect 460 687 461 697
rect 463 687 464 697
rect -1198 665 -1178 666
rect -1198 662 -1178 663
rect -1092 665 -1072 666
rect -1198 657 -1178 658
rect -1326 641 -1325 651
rect -1323 641 -1322 651
rect -1275 641 -1274 651
rect -1272 641 -1271 651
rect -1198 654 -1178 655
rect -1092 662 -1072 663
rect -1092 657 -1072 658
rect -1092 654 -1072 655
rect -871 665 -851 666
rect -871 662 -851 663
rect -765 665 -745 666
rect -871 657 -851 658
rect -998 641 -997 651
rect -995 641 -994 651
rect -948 641 -947 651
rect -945 641 -944 651
rect -871 654 -851 655
rect -765 662 -745 663
rect -765 657 -745 658
rect -765 654 -745 655
rect -539 664 -519 665
rect -539 661 -519 662
rect -433 664 -413 665
rect -539 656 -519 657
rect -667 640 -666 650
rect -664 640 -663 650
rect -616 640 -615 650
rect -613 640 -612 650
rect -539 653 -519 654
rect -433 661 -413 662
rect -433 656 -413 657
rect -433 653 -413 654
rect -212 664 -192 665
rect -212 661 -192 662
rect -106 664 -86 665
rect -212 656 -192 657
rect -339 640 -338 650
rect -336 640 -335 650
rect -289 640 -288 650
rect -286 640 -285 650
rect -212 653 -192 654
rect -106 661 -86 662
rect -106 656 -86 657
rect -106 653 -86 654
rect 691 672 711 673
rect 691 669 711 670
rect 691 664 711 665
rect 691 661 711 662
rect 91 645 111 646
rect 91 642 111 643
rect 91 637 111 638
rect 91 634 111 635
rect 135 625 136 635
rect 138 625 139 635
rect 600 638 620 639
rect 332 632 352 633
rect 332 629 352 630
rect 600 635 620 636
rect 787 638 807 639
rect 600 630 620 631
rect 332 624 352 625
rect 600 627 620 628
rect 787 635 807 636
rect 787 630 807 631
rect 787 627 807 628
rect 332 621 352 622
rect 691 616 711 617
rect 691 613 711 614
rect 691 608 711 609
rect 241 598 261 599
rect 241 595 261 596
rect 691 605 711 606
rect 428 598 448 599
rect 241 590 261 591
rect 241 587 261 588
rect 428 595 448 596
rect 428 590 448 591
rect 428 587 448 588
rect 332 576 352 577
rect 332 573 352 574
rect 332 568 352 569
rect 332 565 352 566
rect 581 534 601 535
rect 581 531 601 532
rect 581 526 601 527
rect -1092 516 -1072 517
rect -1092 513 -1072 514
rect -765 516 -745 517
rect -1092 508 -1072 509
rect -1092 505 -1072 506
rect -765 513 -745 514
rect -433 515 -413 516
rect -765 508 -745 509
rect -1198 498 -1178 499
rect -1198 495 -1178 496
rect -765 505 -745 506
rect -433 512 -413 513
rect 581 523 601 524
rect -106 515 -86 516
rect 625 514 626 524
rect 628 514 629 524
rect -433 507 -413 508
rect -871 498 -851 499
rect -1198 490 -1178 491
rect -1198 487 -1178 488
rect -871 495 -851 496
rect -433 504 -413 505
rect -106 512 -86 513
rect -106 507 -86 508
rect -539 497 -519 498
rect -871 490 -851 491
rect -871 487 -851 488
rect -539 494 -519 495
rect -106 504 -86 505
rect 200 505 220 506
rect -212 497 -192 498
rect -539 489 -519 490
rect -539 486 -519 487
rect -212 494 -192 495
rect 200 502 220 503
rect 200 497 220 498
rect 200 494 220 495
rect -212 489 -192 490
rect -212 486 -192 487
rect 411 483 451 484
rect -1198 451 -1178 452
rect -1198 448 -1178 449
rect -1092 451 -1072 452
rect -1198 443 -1178 444
rect -1326 427 -1325 437
rect -1323 427 -1322 437
rect -1275 427 -1274 437
rect -1272 427 -1271 437
rect -1198 440 -1178 441
rect -1092 448 -1072 449
rect -1092 443 -1072 444
rect -1092 440 -1072 441
rect -871 451 -851 452
rect -871 448 -851 449
rect -765 451 -745 452
rect -871 443 -851 444
rect -998 427 -997 437
rect -995 427 -994 437
rect -948 427 -947 437
rect -945 427 -944 437
rect -871 440 -851 441
rect -765 448 -745 449
rect -765 443 -745 444
rect -765 440 -745 441
rect -539 450 -519 451
rect -539 447 -519 448
rect -433 450 -413 451
rect 109 471 129 472
rect 109 468 129 469
rect 411 480 451 481
rect 411 475 451 476
rect 580 481 610 482
rect 296 471 316 472
rect 109 463 129 464
rect 109 460 129 461
rect 296 468 316 469
rect 411 472 451 473
rect 411 467 451 468
rect 296 463 316 464
rect 296 460 316 461
rect 411 464 451 465
rect 411 459 451 460
rect 580 478 610 479
rect 787 497 797 498
rect 787 494 797 495
rect 787 489 797 490
rect 787 486 797 487
rect 787 481 797 482
rect 580 473 610 474
rect 580 470 610 471
rect 580 465 610 466
rect -539 442 -519 443
rect -667 426 -666 436
rect -664 426 -663 436
rect -616 426 -615 436
rect -613 426 -612 436
rect -539 439 -519 440
rect -433 447 -413 448
rect -433 442 -413 443
rect -433 439 -413 440
rect -212 450 -192 451
rect -212 447 -192 448
rect -106 450 -86 451
rect -212 442 -192 443
rect -339 426 -338 436
rect -336 426 -335 436
rect -289 426 -288 436
rect -286 426 -285 436
rect -212 439 -192 440
rect -106 447 -86 448
rect 411 456 451 457
rect 200 449 220 450
rect 475 449 476 459
rect 478 449 479 459
rect 580 462 610 463
rect 787 478 797 479
rect 787 473 797 474
rect 787 470 797 471
rect 822 461 823 471
rect 825 461 826 471
rect 634 450 635 460
rect 637 450 638 460
rect -106 442 -86 443
rect -106 439 -86 440
rect 200 446 220 447
rect 200 441 220 442
rect 200 438 220 439
rect 758 413 778 414
rect 758 410 778 411
rect 758 405 778 406
rect 758 402 778 403
rect 91 391 111 392
rect 91 388 111 389
rect 91 383 111 384
rect 802 393 803 403
rect 805 393 806 403
rect 91 380 111 381
rect 135 371 136 381
rect 138 371 139 381
rect 339 370 364 371
rect 339 367 364 368
rect 475 372 515 373
rect 339 362 364 363
rect 339 359 364 360
rect 339 354 364 355
rect 339 351 364 352
rect 475 369 515 370
rect 475 364 515 365
rect 621 369 651 370
rect 475 361 515 362
rect 475 356 515 357
rect 339 346 364 347
rect 339 343 364 344
rect 339 338 364 339
rect 389 337 390 347
rect 392 337 393 347
rect 475 353 515 354
rect 475 348 515 349
rect 621 366 651 367
rect 621 361 651 362
rect 621 358 651 359
rect 621 353 651 354
rect 475 345 515 346
rect 539 338 540 348
rect 542 338 543 348
rect 621 350 651 351
rect 675 338 676 348
rect 678 338 679 348
rect 847 349 857 350
rect 847 346 857 347
rect 847 341 857 342
rect 339 335 364 336
rect 847 338 857 339
rect 847 333 857 334
rect 201 323 221 324
rect 847 330 857 331
rect 847 325 857 326
rect 201 320 221 321
rect 201 315 221 316
rect 847 322 857 323
rect 847 317 857 318
rect 880 317 881 327
rect 883 317 884 327
rect 201 312 221 313
rect 847 314 857 315
rect 110 289 130 290
rect -1092 277 -1072 278
rect -1092 274 -1072 275
rect -765 277 -745 278
rect -1092 269 -1072 270
rect -1092 266 -1072 267
rect -765 274 -745 275
rect -433 276 -413 277
rect -765 269 -745 270
rect -1198 259 -1178 260
rect -1198 256 -1178 257
rect -765 266 -745 267
rect -433 273 -413 274
rect 110 286 130 287
rect 297 289 317 290
rect 110 281 130 282
rect -106 276 -86 277
rect 110 278 130 279
rect 297 286 317 287
rect 297 281 317 282
rect 297 278 317 279
rect -433 268 -413 269
rect -871 259 -851 260
rect -1198 251 -1178 252
rect -1198 248 -1178 249
rect -871 256 -851 257
rect -433 265 -413 266
rect -106 273 -86 274
rect -106 268 -86 269
rect -539 258 -519 259
rect -871 251 -851 252
rect -871 248 -851 249
rect -539 255 -519 256
rect -106 265 -86 266
rect 201 267 221 268
rect -212 258 -192 259
rect 201 264 221 265
rect 201 259 221 260
rect -539 250 -519 251
rect -539 247 -519 248
rect -212 255 -192 256
rect 201 256 221 257
rect 524 254 544 255
rect -212 250 -192 251
rect -212 247 -192 248
rect 524 251 544 252
rect 1149 251 1169 252
rect 524 246 544 247
rect 524 243 544 244
rect 1149 248 1169 249
rect 1149 243 1169 244
rect -1198 212 -1178 213
rect -1198 209 -1178 210
rect -1092 212 -1072 213
rect -1198 204 -1178 205
rect -1326 188 -1325 198
rect -1323 188 -1322 198
rect -1275 188 -1274 198
rect -1272 188 -1271 198
rect -1198 201 -1178 202
rect -1092 209 -1072 210
rect -1092 204 -1072 205
rect -1092 201 -1072 202
rect -871 212 -851 213
rect -871 209 -851 210
rect -765 212 -745 213
rect -871 204 -851 205
rect -998 188 -997 198
rect -995 188 -994 198
rect -948 188 -947 198
rect -945 188 -944 198
rect -871 201 -851 202
rect -765 209 -745 210
rect -765 204 -745 205
rect -765 201 -745 202
rect -539 211 -519 212
rect -539 208 -519 209
rect -433 211 -413 212
rect -539 203 -519 204
rect -667 187 -666 197
rect -664 187 -663 197
rect -616 187 -615 197
rect -613 187 -612 197
rect -539 200 -519 201
rect -433 208 -413 209
rect -433 203 -413 204
rect -433 200 -413 201
rect -212 211 -192 212
rect -212 208 -192 209
rect 433 220 453 221
rect -106 211 -86 212
rect -212 203 -192 204
rect -339 187 -338 197
rect -336 187 -335 197
rect -289 187 -288 197
rect -286 187 -285 197
rect -212 200 -192 201
rect -106 208 -86 209
rect 92 209 112 210
rect -106 203 -86 204
rect -106 200 -86 201
rect 92 206 112 207
rect 92 201 112 202
rect 433 217 453 218
rect 620 220 640 221
rect 1149 240 1169 241
rect 433 212 453 213
rect 433 209 453 210
rect 620 217 640 218
rect 620 212 640 213
rect 620 209 640 210
rect 92 198 112 199
rect 136 189 137 199
rect 139 189 140 199
rect 524 198 544 199
rect 738 201 768 202
rect 524 195 544 196
rect 524 190 544 191
rect 738 198 768 199
rect 885 213 905 214
rect 885 210 905 211
rect 885 205 905 206
rect 1058 217 1078 218
rect 1058 214 1078 215
rect 1245 217 1265 218
rect 1058 209 1078 210
rect 885 202 905 203
rect 738 193 768 194
rect 524 187 544 188
rect 738 190 768 191
rect 738 185 768 186
rect 738 182 768 183
rect 929 193 930 203
rect 932 193 933 203
rect 1058 206 1078 207
rect 1245 214 1265 215
rect 1245 209 1265 210
rect 1245 206 1265 207
rect 1149 195 1169 196
rect 1149 192 1169 193
rect 1149 187 1169 188
rect 1149 184 1169 185
rect 792 170 793 180
rect 795 170 796 180
rect 202 140 222 141
rect 202 137 222 138
rect 202 132 222 133
rect 202 129 222 130
rect 413 130 443 131
rect 413 127 443 128
rect 413 122 443 123
rect 413 119 443 120
rect 557 132 582 133
rect 557 129 582 130
rect 557 124 582 125
rect 413 114 443 115
rect 111 106 131 107
rect 111 103 131 104
rect 298 106 318 107
rect 111 98 131 99
rect -1092 90 -1072 91
rect -1092 87 -1072 88
rect -765 90 -745 91
rect -1092 82 -1072 83
rect -1092 79 -1072 80
rect -765 87 -745 88
rect -433 89 -413 90
rect -765 82 -745 83
rect -1198 72 -1178 73
rect -1198 69 -1178 70
rect -765 79 -745 80
rect -433 86 -413 87
rect 111 95 131 96
rect 298 103 318 104
rect 413 111 443 112
rect 413 106 443 107
rect 298 98 318 99
rect 298 95 318 96
rect 413 103 443 104
rect 557 121 582 122
rect 557 116 582 117
rect 557 113 582 114
rect 685 124 725 125
rect 685 121 725 122
rect 685 116 725 117
rect 996 128 1006 129
rect 996 125 1006 126
rect 996 120 1006 121
rect 557 108 582 109
rect 413 98 443 99
rect -106 89 -86 90
rect -433 81 -413 82
rect -871 72 -851 73
rect -1198 64 -1178 65
rect -1198 61 -1178 62
rect -871 69 -851 70
rect -433 78 -413 79
rect -106 86 -86 87
rect -106 81 -86 82
rect 413 95 443 96
rect 413 90 443 91
rect 474 90 475 100
rect 477 90 478 100
rect 557 105 582 106
rect 557 100 582 101
rect 607 99 608 109
rect 610 99 611 109
rect 685 113 725 114
rect 685 108 725 109
rect 557 97 582 98
rect 685 105 725 106
rect 685 100 725 101
rect 996 117 1006 118
rect 996 112 1006 113
rect 996 109 1006 110
rect 996 104 1006 105
rect 685 97 725 98
rect 749 90 750 100
rect 752 90 753 100
rect 996 101 1006 102
rect 996 96 1006 97
rect 202 84 222 85
rect 413 87 443 88
rect 996 93 1006 94
rect 996 88 1006 89
rect 1038 88 1039 98
rect 1041 88 1042 98
rect -539 71 -519 72
rect -871 64 -851 65
rect -871 61 -851 62
rect -539 68 -519 69
rect -106 78 -86 79
rect 202 81 222 82
rect 996 85 1006 86
rect 202 76 222 77
rect -212 71 -192 72
rect 202 73 222 74
rect -539 63 -519 64
rect -539 60 -519 61
rect -212 68 -192 69
rect -212 63 -192 64
rect -212 60 -192 61
rect -1198 25 -1178 26
rect -1198 22 -1178 23
rect -1092 25 -1072 26
rect -1198 17 -1178 18
rect -1326 1 -1325 11
rect -1323 1 -1322 11
rect -1275 1 -1274 11
rect -1272 1 -1271 11
rect -1198 14 -1178 15
rect -1092 22 -1072 23
rect -1092 17 -1072 18
rect -1092 14 -1072 15
rect -871 25 -851 26
rect -871 22 -851 23
rect -765 25 -745 26
rect -871 17 -851 18
rect -998 1 -997 11
rect -995 1 -994 11
rect -948 1 -947 11
rect -945 1 -944 11
rect -871 14 -851 15
rect -765 22 -745 23
rect -765 17 -745 18
rect -765 14 -745 15
rect -539 24 -519 25
rect -539 21 -519 22
rect -433 24 -413 25
rect -539 16 -519 17
rect -667 0 -666 10
rect -664 0 -663 10
rect -616 0 -615 10
rect -613 0 -612 10
rect -539 13 -519 14
rect -433 21 -413 22
rect -433 16 -413 17
rect -433 13 -413 14
rect -212 24 -192 25
rect -212 21 -192 22
rect -106 24 -86 25
rect 93 26 113 27
rect -212 16 -192 17
rect -339 0 -338 10
rect -336 0 -335 10
rect -289 0 -288 10
rect -286 0 -285 10
rect -212 13 -192 14
rect -106 21 -86 22
rect -106 16 -86 17
rect 93 23 113 24
rect 93 18 113 19
rect -106 13 -86 14
rect 93 15 113 16
rect 137 6 138 16
rect 140 6 141 16
<< pdiffusion >>
rect 659 1277 660 1297
rect 662 1277 663 1297
rect 667 1277 668 1297
rect 670 1277 671 1297
rect 724 1277 725 1297
rect 727 1277 728 1297
rect 732 1277 733 1297
rect 735 1277 736 1297
rect 801 1277 802 1297
rect 804 1277 805 1297
rect 809 1277 810 1297
rect 812 1277 813 1297
rect 866 1277 867 1297
rect 869 1277 870 1297
rect 874 1277 875 1297
rect 877 1277 878 1297
rect 941 1277 942 1297
rect 944 1277 945 1297
rect 949 1277 950 1297
rect 952 1277 953 1297
rect 1006 1277 1007 1297
rect 1009 1277 1010 1297
rect 1014 1277 1015 1297
rect 1017 1277 1018 1297
rect 1086 1277 1087 1297
rect 1089 1277 1090 1297
rect 1094 1277 1095 1297
rect 1097 1277 1098 1297
rect 1151 1277 1152 1297
rect 1154 1277 1155 1297
rect 1159 1277 1160 1297
rect 1162 1277 1163 1297
rect 1231 1277 1232 1297
rect 1234 1277 1235 1297
rect 1239 1277 1240 1297
rect 1242 1277 1243 1297
rect 1296 1277 1297 1297
rect 1299 1277 1300 1297
rect 1304 1277 1305 1297
rect 1307 1277 1308 1297
rect 1376 1277 1377 1297
rect 1379 1277 1380 1297
rect 1384 1277 1385 1297
rect 1387 1277 1388 1297
rect 1441 1277 1442 1297
rect 1444 1277 1445 1297
rect 1449 1277 1450 1297
rect 1452 1277 1453 1297
rect 677 1171 678 1191
rect 680 1171 681 1191
rect 685 1171 686 1191
rect 688 1171 689 1191
rect 724 1171 725 1191
rect 727 1171 728 1191
rect 732 1171 733 1191
rect 735 1171 736 1191
rect 819 1171 820 1191
rect 822 1171 823 1191
rect 827 1171 828 1191
rect 830 1171 831 1191
rect 866 1171 867 1191
rect 869 1171 870 1191
rect 874 1171 875 1191
rect 877 1171 878 1191
rect 959 1171 960 1191
rect 962 1171 963 1191
rect 967 1171 968 1191
rect 970 1171 971 1191
rect 1006 1171 1007 1191
rect 1009 1171 1010 1191
rect 1014 1171 1015 1191
rect 1017 1171 1018 1191
rect 1104 1171 1105 1191
rect 1107 1171 1108 1191
rect 1112 1171 1113 1191
rect 1115 1171 1116 1191
rect 1151 1171 1152 1191
rect 1154 1171 1155 1191
rect 1159 1171 1160 1191
rect 1162 1171 1163 1191
rect 1249 1171 1250 1191
rect 1252 1171 1253 1191
rect 1257 1171 1258 1191
rect 1260 1171 1261 1191
rect 1296 1171 1297 1191
rect 1299 1171 1300 1191
rect 1304 1171 1305 1191
rect 1307 1171 1308 1191
rect 1394 1171 1395 1191
rect 1397 1171 1398 1191
rect 1402 1171 1403 1191
rect 1405 1171 1406 1191
rect 1441 1171 1442 1191
rect 1444 1171 1445 1191
rect 1449 1171 1450 1191
rect 1452 1171 1453 1191
rect -468 1129 -448 1130
rect -468 1126 -448 1127
rect -468 1121 -448 1122
rect -141 1129 -121 1130
rect 705 1133 725 1134
rect 847 1133 867 1134
rect 987 1133 1007 1134
rect 1132 1133 1152 1134
rect 1277 1133 1297 1134
rect 1422 1133 1442 1134
rect 705 1130 725 1131
rect -141 1126 -121 1127
rect -468 1118 -448 1119
rect -574 1111 -554 1112
rect -141 1121 -121 1122
rect 847 1130 867 1131
rect 987 1130 1007 1131
rect 1132 1130 1152 1131
rect 1277 1130 1297 1131
rect 1422 1130 1442 1131
rect -141 1118 -121 1119
rect -574 1108 -554 1109
rect -574 1103 -554 1104
rect -247 1111 -227 1112
rect -247 1108 -227 1109
rect -574 1100 -554 1101
rect -247 1103 -227 1104
rect -247 1100 -227 1101
rect -666 1064 -665 1084
rect -663 1064 -662 1084
rect -615 1064 -614 1084
rect -612 1064 -611 1084
rect -574 1064 -554 1065
rect -574 1061 -554 1062
rect -574 1056 -554 1057
rect -468 1064 -448 1065
rect -338 1064 -337 1084
rect -335 1064 -334 1084
rect -288 1064 -287 1084
rect -285 1064 -284 1084
rect 705 1083 725 1084
rect 847 1083 867 1084
rect 987 1083 1007 1084
rect 1132 1083 1152 1084
rect 1277 1083 1297 1084
rect 1422 1083 1442 1084
rect 705 1080 725 1081
rect 847 1080 867 1081
rect 987 1080 1007 1081
rect 1132 1080 1152 1081
rect 1277 1080 1297 1081
rect 1422 1080 1442 1081
rect -468 1061 -448 1062
rect -574 1053 -554 1054
rect -468 1056 -448 1057
rect -468 1053 -448 1054
rect -247 1064 -227 1065
rect -247 1061 -227 1062
rect -247 1056 -227 1057
rect -141 1064 -121 1065
rect -141 1061 -121 1062
rect -247 1053 -227 1054
rect -141 1056 -121 1057
rect -141 1053 -121 1054
rect 416 1027 436 1028
rect 416 1024 436 1025
rect 416 1019 436 1020
rect 416 1016 436 1017
rect 325 993 345 994
rect 325 990 345 991
rect 325 985 345 986
rect 512 993 532 994
rect 512 990 532 991
rect 325 982 345 983
rect 512 985 532 986
rect 512 982 532 983
rect -1128 969 -1108 970
rect -1128 966 -1108 967
rect -1128 961 -1108 962
rect -801 969 -781 970
rect -801 966 -781 967
rect -1128 958 -1108 959
rect -1234 951 -1214 952
rect -801 961 -781 962
rect -469 965 -449 966
rect -469 962 -449 963
rect -801 958 -781 959
rect -1234 948 -1214 949
rect -1234 943 -1214 944
rect -907 951 -887 952
rect -469 957 -449 958
rect -142 965 -122 966
rect 416 971 436 972
rect 416 968 436 969
rect -142 962 -122 963
rect -469 954 -449 955
rect -907 948 -887 949
rect -1234 940 -1214 941
rect -907 943 -887 944
rect -575 947 -555 948
rect -142 957 -122 958
rect 416 963 436 964
rect 416 960 436 961
rect -142 954 -122 955
rect -575 944 -555 945
rect -907 940 -887 941
rect -575 939 -555 940
rect -248 947 -228 948
rect 659 950 660 970
rect 662 950 663 970
rect 667 950 668 970
rect 670 950 671 970
rect 724 950 725 970
rect 727 950 728 970
rect 732 950 733 970
rect 735 950 736 970
rect 801 950 802 970
rect 804 950 805 970
rect 809 950 810 970
rect 812 950 813 970
rect 866 950 867 970
rect 869 950 870 970
rect 874 950 875 970
rect 877 950 878 970
rect 941 950 942 970
rect 944 950 945 970
rect 949 950 950 970
rect 952 950 953 970
rect 1006 950 1007 970
rect 1009 950 1010 970
rect 1014 950 1015 970
rect 1017 950 1018 970
rect 1086 950 1087 970
rect 1089 950 1090 970
rect 1094 950 1095 970
rect 1097 950 1098 970
rect 1151 950 1152 970
rect 1154 950 1155 970
rect 1159 950 1160 970
rect 1162 950 1163 970
rect 1231 950 1232 970
rect 1234 950 1235 970
rect 1239 950 1240 970
rect 1242 950 1243 970
rect 1296 950 1297 970
rect 1299 950 1300 970
rect 1304 950 1305 970
rect 1307 950 1308 970
rect 1376 950 1377 970
rect 1379 950 1380 970
rect 1384 950 1385 970
rect 1387 950 1388 970
rect 1441 950 1442 970
rect 1444 950 1445 970
rect 1449 950 1450 970
rect 1452 950 1453 970
rect -248 944 -228 945
rect -575 936 -555 937
rect -248 939 -228 940
rect -248 936 -228 937
rect 165 939 185 940
rect 165 936 185 937
rect 165 931 185 932
rect 165 928 185 929
rect -1326 904 -1325 924
rect -1323 904 -1322 924
rect -1275 904 -1274 924
rect -1272 904 -1271 924
rect -1234 904 -1214 905
rect -1234 901 -1214 902
rect -1234 896 -1214 897
rect -1128 904 -1108 905
rect -998 904 -997 924
rect -995 904 -994 924
rect -948 904 -947 924
rect -945 904 -944 924
rect -1128 901 -1108 902
rect -1234 893 -1214 894
rect -1128 896 -1108 897
rect -1128 893 -1108 894
rect -907 904 -887 905
rect -907 901 -887 902
rect -907 896 -887 897
rect -801 904 -781 905
rect -801 901 -781 902
rect -907 893 -887 894
rect -801 896 -781 897
rect -667 900 -666 920
rect -664 900 -663 920
rect -616 900 -615 920
rect -613 900 -612 920
rect -801 893 -781 894
rect -575 900 -555 901
rect -575 897 -555 898
rect -575 892 -555 893
rect -469 900 -449 901
rect -339 900 -338 920
rect -336 900 -335 920
rect -289 900 -288 920
rect -286 900 -285 920
rect -469 897 -449 898
rect -575 889 -555 890
rect -469 892 -449 893
rect -469 889 -449 890
rect -248 900 -228 901
rect -248 897 -228 898
rect -248 892 -228 893
rect -142 900 -122 901
rect 74 905 94 906
rect 74 902 94 903
rect -142 897 -122 898
rect -248 889 -228 890
rect -142 892 -122 893
rect 74 897 94 898
rect 261 905 281 906
rect 261 902 281 903
rect 74 894 94 895
rect 261 897 281 898
rect 261 894 281 895
rect 445 892 446 912
rect 448 892 449 912
rect 573 892 574 912
rect 576 892 577 912
rect -142 889 -122 890
rect 165 883 185 884
rect 368 886 388 887
rect 368 883 388 884
rect 165 880 185 881
rect 165 875 185 876
rect 368 878 388 879
rect 486 885 526 886
rect 486 882 526 883
rect 368 875 388 876
rect 165 872 185 873
rect 486 877 526 878
rect 486 874 526 875
rect 136 831 137 851
rect 139 831 140 851
rect 677 844 678 864
rect 680 844 681 864
rect 685 844 686 864
rect 688 844 689 864
rect 724 844 725 864
rect 727 844 728 864
rect 732 844 733 864
rect 735 844 736 864
rect 819 844 820 864
rect 822 844 823 864
rect 827 844 828 864
rect 830 844 831 864
rect 866 844 867 864
rect 869 844 870 864
rect 874 844 875 864
rect 877 844 878 864
rect 959 844 960 864
rect 962 844 963 864
rect 967 844 968 864
rect 970 844 971 864
rect 1006 844 1007 864
rect 1009 844 1010 864
rect 1014 844 1015 864
rect 1017 844 1018 864
rect 1104 844 1105 864
rect 1107 844 1108 864
rect 1112 844 1113 864
rect 1115 844 1116 864
rect 1151 844 1152 864
rect 1154 844 1155 864
rect 1159 844 1160 864
rect 1162 844 1163 864
rect 1249 844 1250 864
rect 1252 844 1253 864
rect 1257 844 1258 864
rect 1260 844 1261 864
rect 1296 844 1297 864
rect 1299 844 1300 864
rect 1304 844 1305 864
rect 1307 844 1308 864
rect 1394 844 1395 864
rect 1397 844 1398 864
rect 1402 844 1403 864
rect 1405 844 1406 864
rect 1441 844 1442 864
rect 1444 844 1445 864
rect 1449 844 1450 864
rect 1452 844 1453 864
rect 59 825 79 826
rect 59 822 79 823
rect 59 817 79 818
rect 59 814 79 815
rect 368 806 369 826
rect 371 806 372 826
rect 291 800 311 801
rect 291 797 311 798
rect 291 792 311 793
rect 415 803 475 804
rect 415 800 475 801
rect 415 795 475 796
rect 521 799 522 819
rect 524 799 525 819
rect 705 806 725 807
rect 847 806 867 807
rect 987 806 1007 807
rect 1132 806 1152 807
rect 1277 806 1297 807
rect 1422 806 1442 807
rect 705 803 725 804
rect 847 803 867 804
rect 987 803 1007 804
rect 1132 803 1152 804
rect 1277 803 1297 804
rect 1422 803 1442 804
rect 415 792 475 793
rect 291 789 311 790
rect 415 787 475 788
rect 415 784 475 785
rect 164 759 184 760
rect 164 756 184 757
rect 164 751 184 752
rect 705 755 725 756
rect 847 755 867 756
rect 987 755 1007 756
rect 1132 755 1152 756
rect 1277 755 1297 756
rect 1422 755 1442 756
rect 705 752 725 753
rect 164 748 184 749
rect 847 752 867 753
rect 987 752 1007 753
rect 1132 752 1152 753
rect 1277 752 1297 753
rect 1422 752 1442 753
rect -1128 730 -1108 731
rect -1128 727 -1108 728
rect -1128 722 -1108 723
rect -801 730 -781 731
rect -801 727 -781 728
rect -1128 719 -1108 720
rect -1234 712 -1214 713
rect -801 722 -781 723
rect -469 729 -449 730
rect -469 726 -449 727
rect -801 719 -781 720
rect -1234 709 -1214 710
rect -1234 704 -1214 705
rect -907 712 -887 713
rect -469 721 -449 722
rect -142 729 -122 730
rect -142 726 -122 727
rect -469 718 -449 719
rect -907 709 -887 710
rect -1234 701 -1214 702
rect -907 704 -887 705
rect -575 711 -555 712
rect -142 721 -122 722
rect 73 725 93 726
rect 73 722 93 723
rect -142 718 -122 719
rect -575 708 -555 709
rect -907 701 -887 702
rect -575 703 -555 704
rect -248 711 -228 712
rect 73 717 93 718
rect 260 725 280 726
rect 260 722 280 723
rect 73 714 93 715
rect 260 717 280 718
rect 374 718 394 719
rect 374 715 394 716
rect 260 714 280 715
rect -248 708 -228 709
rect -575 700 -555 701
rect -248 703 -228 704
rect -248 700 -228 701
rect 164 703 184 704
rect 374 710 394 711
rect 460 713 461 733
rect 463 713 464 733
rect 374 707 394 708
rect 164 700 184 701
rect 164 695 184 696
rect 374 702 394 703
rect 374 699 394 700
rect 164 692 184 693
rect -1326 665 -1325 685
rect -1323 665 -1322 685
rect -1275 665 -1274 685
rect -1272 665 -1271 685
rect -1234 665 -1214 666
rect -1234 662 -1214 663
rect -1234 657 -1214 658
rect -1128 665 -1108 666
rect -998 665 -997 685
rect -995 665 -994 685
rect -948 665 -947 685
rect -945 665 -944 685
rect -1128 662 -1108 663
rect -1234 654 -1214 655
rect -1128 657 -1108 658
rect -1128 654 -1108 655
rect -907 665 -887 666
rect -907 662 -887 663
rect -907 657 -887 658
rect -801 665 -781 666
rect -667 664 -666 684
rect -664 664 -663 684
rect -616 664 -615 684
rect -613 664 -612 684
rect -801 662 -781 663
rect -907 654 -887 655
rect -801 657 -781 658
rect -801 654 -781 655
rect -575 664 -555 665
rect -575 661 -555 662
rect -575 656 -555 657
rect -469 664 -449 665
rect -339 664 -338 684
rect -336 664 -335 684
rect -289 664 -288 684
rect -286 664 -285 684
rect -469 661 -449 662
rect -575 653 -555 654
rect -469 656 -449 657
rect -469 653 -449 654
rect -248 664 -228 665
rect -248 661 -228 662
rect -248 656 -228 657
rect -142 664 -122 665
rect -142 661 -122 662
rect -248 653 -228 654
rect -142 656 -122 657
rect -142 653 -122 654
rect 135 651 136 671
rect 138 651 139 671
rect 655 672 675 673
rect 655 669 675 670
rect 655 664 675 665
rect 655 661 675 662
rect 58 645 78 646
rect 58 642 78 643
rect 58 637 78 638
rect 58 634 78 635
rect 296 632 316 633
rect 564 638 584 639
rect 564 635 584 636
rect 296 629 316 630
rect 296 624 316 625
rect 564 630 584 631
rect 751 638 771 639
rect 751 635 771 636
rect 564 627 584 628
rect 751 630 771 631
rect 751 627 771 628
rect 296 621 316 622
rect 655 616 675 617
rect 655 613 675 614
rect 655 608 675 609
rect 655 605 675 606
rect 205 598 225 599
rect 205 595 225 596
rect 205 590 225 591
rect 392 598 412 599
rect 392 595 412 596
rect 205 587 225 588
rect 392 590 412 591
rect 392 587 412 588
rect 296 576 316 577
rect 296 573 316 574
rect 296 568 316 569
rect 296 565 316 566
rect 625 540 626 560
rect 628 540 629 560
rect 548 534 568 535
rect 548 531 568 532
rect 548 526 568 527
rect 548 523 568 524
rect -1128 516 -1108 517
rect -1128 513 -1108 514
rect -1128 508 -1108 509
rect -801 516 -781 517
rect -801 513 -781 514
rect -1128 505 -1108 506
rect -1234 498 -1214 499
rect -801 508 -781 509
rect -469 515 -449 516
rect -469 512 -449 513
rect -801 505 -781 506
rect -1234 495 -1214 496
rect -1234 490 -1214 491
rect -907 498 -887 499
rect -469 507 -449 508
rect -142 515 -122 516
rect -142 512 -122 513
rect -469 504 -449 505
rect -907 495 -887 496
rect -1234 487 -1214 488
rect -907 490 -887 491
rect -575 497 -555 498
rect -142 507 -122 508
rect -142 504 -122 505
rect -575 494 -555 495
rect -907 487 -887 488
rect -575 489 -555 490
rect -248 497 -228 498
rect 164 505 184 506
rect 164 502 184 503
rect -248 494 -228 495
rect -575 486 -555 487
rect -248 489 -228 490
rect 164 497 184 498
rect 164 494 184 495
rect -248 486 -228 487
rect 379 483 399 484
rect 379 480 399 481
rect -1326 451 -1325 471
rect -1323 451 -1322 471
rect -1275 451 -1274 471
rect -1272 451 -1271 471
rect -1234 451 -1214 452
rect -1234 448 -1214 449
rect -1234 443 -1214 444
rect -1128 451 -1108 452
rect -998 451 -997 471
rect -995 451 -994 471
rect -948 451 -947 471
rect -945 451 -944 471
rect -1128 448 -1108 449
rect -1234 440 -1214 441
rect -1128 443 -1108 444
rect -1128 440 -1108 441
rect -907 451 -887 452
rect -907 448 -887 449
rect -907 443 -887 444
rect -801 451 -781 452
rect -667 450 -666 470
rect -664 450 -663 470
rect -616 450 -615 470
rect -613 450 -612 470
rect -801 448 -781 449
rect -907 440 -887 441
rect -801 443 -781 444
rect -801 440 -781 441
rect -575 450 -555 451
rect -575 447 -555 448
rect -575 442 -555 443
rect -469 450 -449 451
rect -339 450 -338 470
rect -336 450 -335 470
rect -289 450 -288 470
rect -286 450 -285 470
rect 73 471 93 472
rect 73 468 93 469
rect 73 463 93 464
rect 260 471 280 472
rect 379 475 399 476
rect 475 475 476 495
rect 478 475 479 495
rect 548 481 568 482
rect 548 478 568 479
rect 379 472 399 473
rect 260 468 280 469
rect 73 460 93 461
rect 260 463 280 464
rect 379 467 399 468
rect 379 464 399 465
rect 260 460 280 461
rect 379 459 399 460
rect 548 473 568 474
rect 634 476 635 496
rect 637 476 638 496
rect 695 497 775 498
rect 695 494 775 495
rect 695 489 775 490
rect 822 487 823 507
rect 825 487 826 507
rect 695 486 775 487
rect 695 481 775 482
rect 695 478 775 479
rect 548 470 568 471
rect 548 465 568 466
rect 548 462 568 463
rect 379 456 399 457
rect -469 447 -449 448
rect -575 439 -555 440
rect -469 442 -449 443
rect -469 439 -449 440
rect -248 450 -228 451
rect -248 447 -228 448
rect -248 442 -228 443
rect -142 450 -122 451
rect -142 447 -122 448
rect -248 439 -228 440
rect -142 442 -122 443
rect 164 449 184 450
rect 695 473 775 474
rect 695 470 775 471
rect 164 446 184 447
rect -142 439 -122 440
rect 164 441 184 442
rect 164 438 184 439
rect 802 419 803 439
rect 805 419 806 439
rect 135 397 136 417
rect 138 397 139 417
rect 725 413 745 414
rect 725 410 745 411
rect 725 405 745 406
rect 725 402 745 403
rect 58 391 78 392
rect 58 388 78 389
rect 58 383 78 384
rect 58 380 78 381
rect 307 370 327 371
rect 307 367 327 368
rect 307 362 327 363
rect 389 363 390 383
rect 392 363 393 383
rect 443 372 463 373
rect 443 369 463 370
rect 307 359 327 360
rect 307 354 327 355
rect 307 351 327 352
rect 307 346 327 347
rect 443 364 463 365
rect 539 364 540 384
rect 542 364 543 384
rect 589 369 609 370
rect 589 366 609 367
rect 443 361 463 362
rect 443 356 463 357
rect 443 353 463 354
rect 307 343 327 344
rect 307 338 327 339
rect 443 348 463 349
rect 589 361 609 362
rect 675 364 676 384
rect 678 364 679 384
rect 589 358 609 359
rect 589 353 609 354
rect 589 350 609 351
rect 443 345 463 346
rect 735 349 835 350
rect 735 346 835 347
rect 735 341 835 342
rect 880 343 881 363
rect 883 343 884 363
rect 735 338 835 339
rect 307 335 327 336
rect 735 333 835 334
rect 735 330 835 331
rect 165 323 185 324
rect 735 325 835 326
rect 735 322 835 323
rect 165 320 185 321
rect 165 315 185 316
rect 735 317 835 318
rect 735 314 835 315
rect 165 312 185 313
rect 74 289 94 290
rect 74 286 94 287
rect -1128 277 -1108 278
rect -1128 274 -1108 275
rect -1128 269 -1108 270
rect -801 277 -781 278
rect -801 274 -781 275
rect -1128 266 -1108 267
rect -1234 259 -1214 260
rect -801 269 -781 270
rect -469 276 -449 277
rect -469 273 -449 274
rect -801 266 -781 267
rect -1234 256 -1214 257
rect -1234 251 -1214 252
rect -907 259 -887 260
rect -469 268 -449 269
rect -142 276 -122 277
rect 74 281 94 282
rect 261 289 281 290
rect 261 286 281 287
rect 74 278 94 279
rect 261 281 281 282
rect 261 278 281 279
rect -142 273 -122 274
rect -469 265 -449 266
rect -907 256 -887 257
rect -1234 248 -1214 249
rect -907 251 -887 252
rect -575 258 -555 259
rect -142 268 -122 269
rect -142 265 -122 266
rect -575 255 -555 256
rect -907 248 -887 249
rect -575 250 -555 251
rect -248 258 -228 259
rect 165 267 185 268
rect 165 264 185 265
rect 165 259 185 260
rect 165 256 185 257
rect -248 255 -228 256
rect -575 247 -555 248
rect -248 250 -228 251
rect 488 254 508 255
rect 488 251 508 252
rect -248 247 -228 248
rect 488 246 508 247
rect 1113 251 1133 252
rect 1113 248 1133 249
rect 488 243 508 244
rect 1113 243 1133 244
rect 1113 240 1133 241
rect -1326 212 -1325 232
rect -1323 212 -1322 232
rect -1275 212 -1274 232
rect -1272 212 -1271 232
rect -1234 212 -1214 213
rect -1234 209 -1214 210
rect -1234 204 -1214 205
rect -1128 212 -1108 213
rect -998 212 -997 232
rect -995 212 -994 232
rect -948 212 -947 232
rect -945 212 -944 232
rect -1128 209 -1108 210
rect -1234 201 -1214 202
rect -1128 204 -1108 205
rect -1128 201 -1108 202
rect -907 212 -887 213
rect -907 209 -887 210
rect -907 204 -887 205
rect -801 212 -781 213
rect -667 211 -666 231
rect -664 211 -663 231
rect -616 211 -615 231
rect -613 211 -612 231
rect -801 209 -781 210
rect -907 201 -887 202
rect -801 204 -781 205
rect -801 201 -781 202
rect -575 211 -555 212
rect -575 208 -555 209
rect -575 203 -555 204
rect -469 211 -449 212
rect -339 211 -338 231
rect -336 211 -335 231
rect -289 211 -288 231
rect -286 211 -285 231
rect -469 208 -449 209
rect -575 200 -555 201
rect -469 203 -449 204
rect -469 200 -449 201
rect -248 211 -228 212
rect -248 208 -228 209
rect -248 203 -228 204
rect -142 211 -122 212
rect 136 215 137 235
rect 139 215 140 235
rect 397 220 417 221
rect 397 217 417 218
rect -142 208 -122 209
rect -248 200 -228 201
rect -142 203 -122 204
rect 59 209 79 210
rect 59 206 79 207
rect -142 200 -122 201
rect 59 201 79 202
rect 397 212 417 213
rect 584 220 604 221
rect 929 219 930 239
rect 932 219 933 239
rect 584 217 604 218
rect 397 209 417 210
rect 584 212 604 213
rect 584 209 604 210
rect 59 198 79 199
rect 488 198 508 199
rect 706 201 726 202
rect 706 198 726 199
rect 488 195 508 196
rect 488 190 508 191
rect 706 193 726 194
rect 792 196 793 216
rect 795 196 796 216
rect 852 213 872 214
rect 852 210 872 211
rect 852 205 872 206
rect 1022 217 1042 218
rect 1022 214 1042 215
rect 1022 209 1042 210
rect 1209 217 1229 218
rect 1209 214 1229 215
rect 1022 206 1042 207
rect 852 202 872 203
rect 706 190 726 191
rect 488 187 508 188
rect 706 185 726 186
rect 706 182 726 183
rect 1209 209 1229 210
rect 1209 206 1229 207
rect 1113 195 1133 196
rect 1113 192 1133 193
rect 1113 187 1133 188
rect 1113 184 1133 185
rect 166 140 186 141
rect 166 137 186 138
rect 166 132 186 133
rect 166 129 186 130
rect 389 130 399 131
rect 389 127 399 128
rect 389 122 399 123
rect 389 119 399 120
rect 389 114 399 115
rect 474 116 475 136
rect 477 116 478 136
rect 525 132 545 133
rect 525 129 545 130
rect 525 124 545 125
rect 607 125 608 145
rect 610 125 611 145
rect 525 121 545 122
rect 389 111 399 112
rect 75 106 95 107
rect 75 103 95 104
rect 75 98 95 99
rect 262 106 282 107
rect 262 103 282 104
rect 75 95 95 96
rect -1128 90 -1108 91
rect -1128 87 -1108 88
rect -1128 82 -1108 83
rect -801 90 -781 91
rect -801 87 -781 88
rect -1128 79 -1108 80
rect -1234 72 -1214 73
rect -801 82 -781 83
rect -469 89 -449 90
rect -469 86 -449 87
rect -801 79 -781 80
rect -1234 69 -1214 70
rect -1234 64 -1214 65
rect -907 72 -887 73
rect -469 81 -449 82
rect -142 89 -122 90
rect 262 98 282 99
rect 389 106 399 107
rect 389 103 399 104
rect 262 95 282 96
rect 389 98 399 99
rect 525 116 545 117
rect 525 113 545 114
rect 525 108 545 109
rect 653 124 673 125
rect 653 121 673 122
rect 653 116 673 117
rect 749 116 750 136
rect 752 116 753 136
rect 864 128 984 129
rect 864 125 984 126
rect 864 120 984 121
rect 864 117 984 118
rect 653 113 673 114
rect 525 105 545 106
rect 389 95 399 96
rect -142 86 -122 87
rect -469 78 -449 79
rect -907 69 -887 70
rect -1234 61 -1214 62
rect -907 64 -887 65
rect -575 71 -555 72
rect -142 81 -122 82
rect 166 84 186 85
rect 389 90 399 91
rect 525 100 545 101
rect 653 108 673 109
rect 653 105 673 106
rect 525 97 545 98
rect 653 100 673 101
rect 864 112 984 113
rect 1038 114 1039 134
rect 1041 114 1042 134
rect 864 109 984 110
rect 864 104 984 105
rect 864 101 984 102
rect 653 97 673 98
rect 864 96 984 97
rect 864 93 984 94
rect 389 87 399 88
rect 864 88 984 89
rect 864 85 984 86
rect 166 81 186 82
rect -142 78 -122 79
rect -575 68 -555 69
rect -907 61 -887 62
rect -575 63 -555 64
rect -248 71 -228 72
rect 166 76 186 77
rect 166 73 186 74
rect -248 68 -228 69
rect -575 60 -555 61
rect -248 63 -228 64
rect -248 60 -228 61
rect -1326 25 -1325 45
rect -1323 25 -1322 45
rect -1275 25 -1274 45
rect -1272 25 -1271 45
rect -1234 25 -1214 26
rect -1234 22 -1214 23
rect -1234 17 -1214 18
rect -1128 25 -1108 26
rect -998 25 -997 45
rect -995 25 -994 45
rect -948 25 -947 45
rect -945 25 -944 45
rect -1128 22 -1108 23
rect -1234 14 -1214 15
rect -1128 17 -1108 18
rect -1128 14 -1108 15
rect -907 25 -887 26
rect -907 22 -887 23
rect -907 17 -887 18
rect -801 25 -781 26
rect -667 24 -666 44
rect -664 24 -663 44
rect -616 24 -615 44
rect -613 24 -612 44
rect -801 22 -781 23
rect -907 14 -887 15
rect -801 17 -781 18
rect -801 14 -781 15
rect -575 24 -555 25
rect -575 21 -555 22
rect -575 16 -555 17
rect -469 24 -449 25
rect -339 24 -338 44
rect -336 24 -335 44
rect -289 24 -288 44
rect -286 24 -285 44
rect 137 32 138 52
rect 140 32 141 52
rect -469 21 -449 22
rect -575 13 -555 14
rect -469 16 -449 17
rect -469 13 -449 14
rect -248 24 -228 25
rect -248 21 -228 22
rect -248 16 -228 17
rect -142 24 -122 25
rect 60 26 80 27
rect 60 23 80 24
rect -142 21 -122 22
rect -248 13 -228 14
rect -142 16 -122 17
rect 60 18 80 19
rect 60 15 80 16
rect -142 13 -122 14
<< metal1 >>
rect 645 1347 649 1379
rect 659 1353 758 1356
rect 645 1343 690 1347
rect 645 1309 649 1343
rect 655 1333 659 1335
rect 671 1309 675 1313
rect 645 1305 675 1309
rect 663 1297 667 1305
rect 655 1271 659 1277
rect 671 1271 675 1277
rect 641 1268 681 1271
rect 641 1166 644 1268
rect 686 1265 690 1343
rect 720 1333 724 1353
rect 736 1309 740 1313
rect 698 1305 740 1309
rect 728 1297 732 1305
rect 720 1271 724 1277
rect 736 1271 740 1277
rect 714 1268 746 1271
rect 671 1261 678 1264
rect 659 1203 663 1261
rect 686 1261 724 1265
rect 732 1245 736 1261
rect 706 1241 736 1245
rect 667 1233 695 1236
rect 673 1227 677 1233
rect 689 1203 693 1207
rect 659 1199 693 1203
rect 706 1203 710 1241
rect 755 1236 758 1353
rect 787 1347 791 1379
rect 801 1353 900 1356
rect 787 1343 832 1347
rect 787 1309 791 1343
rect 797 1333 801 1335
rect 813 1309 817 1313
rect 787 1305 817 1309
rect 805 1297 809 1305
rect 797 1271 801 1277
rect 813 1271 817 1277
rect 718 1233 758 1236
rect 720 1227 724 1233
rect 736 1203 740 1207
rect 706 1199 740 1203
rect 681 1191 685 1199
rect 728 1191 732 1199
rect 635 1165 644 1166
rect 673 1165 677 1171
rect 689 1165 693 1171
rect 720 1165 724 1171
rect 736 1165 740 1171
rect 635 1162 696 1165
rect -526 1151 -252 1154
rect -526 1148 -523 1151
rect -256 1148 -252 1151
rect -676 1145 -474 1148
rect -583 1116 -580 1145
rect -477 1134 -474 1145
rect -256 1145 -147 1148
rect -440 1140 -304 1144
rect -477 1130 -468 1134
rect -546 1126 -484 1130
rect -583 1112 -574 1116
rect -691 1108 -590 1112
rect -676 1090 -656 1094
rect -670 1084 -666 1090
rect -662 1057 -658 1064
rect -645 1057 -642 1099
rect -691 1053 -669 1057
rect -662 1053 -642 1057
rect -635 1057 -631 1108
rect -620 1090 -606 1094
rect -619 1084 -615 1090
rect -611 1057 -607 1064
rect -594 1061 -590 1104
rect -583 1100 -580 1112
rect -546 1108 -542 1126
rect -512 1116 -509 1122
rect -518 1112 -509 1116
rect -554 1104 -542 1108
rect -546 1100 -542 1104
rect -583 1096 -574 1100
rect -546 1096 -538 1100
rect -583 1093 -580 1096
rect -512 1094 -509 1112
rect -477 1118 -474 1130
rect -440 1126 -436 1140
rect -412 1130 -410 1134
rect -448 1122 -436 1126
rect -440 1118 -436 1122
rect -484 1111 -481 1118
rect -477 1114 -468 1118
rect -440 1114 -432 1118
rect -477 1108 -474 1114
rect -402 1103 -398 1140
rect -484 1099 -398 1103
rect -546 1079 -500 1083
rect -583 1069 -580 1072
rect -583 1065 -574 1069
rect -635 1053 -618 1057
rect -611 1053 -590 1057
rect -583 1053 -580 1065
rect -546 1061 -542 1079
rect -512 1069 -509 1071
rect -518 1065 -509 1069
rect -554 1057 -542 1061
rect -546 1053 -542 1057
rect -662 1050 -658 1053
rect -611 1050 -607 1053
rect -583 1049 -574 1053
rect -546 1049 -538 1053
rect -583 1043 -580 1049
rect -670 1034 -666 1040
rect -619 1034 -615 1040
rect -512 1034 -509 1065
rect -504 1057 -500 1079
rect -484 1065 -480 1099
rect -477 1069 -474 1075
rect -477 1065 -468 1069
rect -504 1053 -484 1057
rect -477 1053 -474 1065
rect -440 1061 -436 1091
rect -392 1069 -389 1130
rect -308 1112 -304 1140
rect -256 1116 -253 1145
rect -150 1134 -147 1145
rect -113 1140 6 1144
rect -150 1130 -141 1134
rect -219 1126 -157 1130
rect -256 1112 -247 1116
rect -308 1108 -263 1112
rect -348 1090 -324 1094
rect -412 1065 -389 1069
rect -448 1057 -436 1061
rect -440 1053 -436 1057
rect -477 1049 -468 1053
rect -440 1049 -432 1053
rect -477 1043 -474 1049
rect -392 1034 -389 1065
rect -342 1084 -338 1090
rect -334 1057 -330 1064
rect -318 1057 -313 1099
rect -353 1053 -341 1057
rect -334 1053 -313 1057
rect -308 1057 -304 1108
rect -293 1090 -279 1094
rect -292 1084 -288 1090
rect -284 1057 -280 1064
rect -267 1061 -263 1104
rect -256 1100 -253 1112
rect -219 1108 -215 1126
rect -185 1116 -182 1122
rect -191 1112 -182 1116
rect -227 1104 -215 1108
rect -219 1100 -215 1104
rect -256 1096 -247 1100
rect -219 1096 -211 1100
rect -256 1093 -253 1096
rect -185 1094 -182 1112
rect -150 1118 -147 1130
rect -113 1126 -109 1140
rect -85 1130 -83 1134
rect -121 1122 -109 1126
rect -113 1118 -109 1122
rect -157 1111 -154 1118
rect -150 1114 -141 1118
rect -113 1114 -105 1118
rect -150 1108 -147 1114
rect -75 1103 -71 1140
rect -157 1099 -71 1103
rect -219 1079 -173 1083
rect -256 1069 -253 1072
rect -256 1065 -247 1069
rect -308 1053 -291 1057
rect -284 1053 -263 1057
rect -256 1053 -253 1065
rect -219 1061 -215 1079
rect -185 1069 -182 1071
rect -191 1065 -182 1069
rect -227 1057 -215 1061
rect -219 1053 -215 1057
rect -334 1050 -330 1053
rect -284 1050 -280 1053
rect -256 1049 -247 1053
rect -219 1049 -211 1053
rect -256 1043 -253 1049
rect -342 1034 -338 1040
rect -292 1034 -288 1040
rect -185 1034 -182 1065
rect -177 1057 -173 1079
rect -157 1065 -153 1099
rect -150 1069 -147 1075
rect -150 1065 -141 1069
rect -177 1053 -157 1057
rect -150 1053 -147 1065
rect -113 1061 -109 1091
rect -65 1069 -62 1130
rect -85 1065 -62 1069
rect -121 1057 -109 1061
rect -113 1053 -109 1057
rect -150 1049 -141 1053
rect -113 1049 -105 1053
rect -150 1043 -147 1049
rect -65 1034 -62 1065
rect -670 1031 -62 1034
rect -703 996 -4 1000
rect -1186 991 -912 994
rect -1186 988 -1183 991
rect -916 988 -912 991
rect -1336 985 -1134 988
rect -1243 956 -1240 985
rect -1137 974 -1134 985
rect -916 985 -807 988
rect -1100 980 -964 984
rect -1137 970 -1128 974
rect -1206 966 -1144 970
rect -1243 952 -1234 956
rect -1351 948 -1250 952
rect -1336 930 -1316 934
rect -1330 924 -1326 930
rect -1322 897 -1318 904
rect -1305 897 -1302 939
rect -1351 893 -1329 897
rect -1322 893 -1302 897
rect -1295 897 -1291 948
rect -1280 930 -1266 934
rect -1279 924 -1275 930
rect -1271 897 -1267 904
rect -1254 901 -1250 944
rect -1243 940 -1240 952
rect -1206 948 -1202 966
rect -1172 956 -1169 962
rect -1178 952 -1169 956
rect -1214 944 -1202 948
rect -1206 940 -1202 944
rect -1243 936 -1234 940
rect -1206 936 -1198 940
rect -1243 933 -1240 936
rect -1172 934 -1169 952
rect -1137 958 -1134 970
rect -1100 966 -1096 980
rect -1072 970 -1070 974
rect -1108 962 -1096 966
rect -1100 958 -1096 962
rect -1144 951 -1141 958
rect -1137 954 -1128 958
rect -1100 954 -1092 958
rect -1137 948 -1134 954
rect -1062 943 -1058 980
rect -1144 939 -1058 943
rect -1206 919 -1160 923
rect -1243 909 -1240 912
rect -1243 905 -1234 909
rect -1295 893 -1278 897
rect -1271 893 -1250 897
rect -1243 893 -1240 905
rect -1206 901 -1202 919
rect -1172 909 -1169 911
rect -1178 905 -1169 909
rect -1214 897 -1202 901
rect -1206 893 -1202 897
rect -1322 890 -1318 893
rect -1271 890 -1267 893
rect -1243 889 -1234 893
rect -1206 889 -1198 893
rect -1243 883 -1240 889
rect -1330 874 -1326 880
rect -1279 874 -1275 880
rect -1172 874 -1169 905
rect -1164 897 -1160 919
rect -1144 905 -1140 939
rect -1137 909 -1134 915
rect -1137 905 -1128 909
rect -1164 893 -1144 897
rect -1137 893 -1134 905
rect -1100 901 -1096 931
rect -1052 909 -1049 970
rect -968 952 -964 980
rect -916 956 -913 985
rect -810 974 -807 985
rect -703 984 -699 996
rect -527 987 -253 990
rect -527 984 -524 987
rect -257 984 -253 987
rect -773 980 -699 984
rect -677 981 -475 984
rect -810 970 -801 974
rect -879 966 -817 970
rect -916 952 -907 956
rect -968 948 -923 952
rect -1008 930 -984 934
rect -1072 905 -1049 909
rect -1108 897 -1096 901
rect -1100 893 -1096 897
rect -1137 889 -1128 893
rect -1100 889 -1092 893
rect -1137 883 -1134 889
rect -1052 874 -1049 905
rect -1002 924 -998 930
rect -994 897 -990 904
rect -978 897 -973 939
rect -1013 893 -1001 897
rect -994 893 -973 897
rect -968 897 -964 948
rect -953 930 -939 934
rect -952 924 -948 930
rect -944 897 -940 904
rect -927 901 -923 944
rect -916 940 -913 952
rect -879 948 -875 966
rect -845 956 -842 962
rect -851 952 -842 956
rect -887 944 -875 948
rect -879 940 -875 944
rect -916 936 -907 940
rect -879 936 -871 940
rect -916 933 -913 936
rect -845 934 -842 952
rect -810 958 -807 970
rect -773 966 -769 980
rect -745 970 -743 974
rect -781 962 -769 966
rect -773 958 -769 962
rect -817 951 -814 958
rect -810 954 -801 958
rect -773 954 -765 958
rect -810 948 -807 954
rect -735 943 -731 980
rect -817 939 -731 943
rect -879 919 -833 923
rect -916 909 -913 912
rect -916 905 -907 909
rect -968 893 -951 897
rect -944 893 -923 897
rect -916 893 -913 905
rect -879 901 -875 919
rect -845 909 -842 911
rect -851 905 -842 909
rect -887 897 -875 901
rect -879 893 -875 897
rect -994 890 -990 893
rect -944 890 -940 893
rect -916 889 -907 893
rect -879 889 -871 893
rect -916 883 -913 889
rect -1002 874 -998 880
rect -952 874 -948 880
rect -845 874 -842 905
rect -837 897 -833 919
rect -817 905 -813 939
rect -810 909 -807 915
rect -810 905 -801 909
rect -837 893 -817 897
rect -810 893 -807 905
rect -773 901 -769 931
rect -725 909 -722 970
rect -584 952 -581 981
rect -478 970 -475 981
rect -257 981 -148 984
rect -441 976 -305 980
rect -478 966 -469 970
rect -547 962 -485 966
rect -584 948 -575 952
rect -692 944 -591 948
rect -677 926 -657 930
rect -745 905 -722 909
rect -781 897 -769 901
rect -773 893 -769 897
rect -810 889 -801 893
rect -773 889 -765 893
rect -810 883 -807 889
rect -725 874 -722 905
rect -671 920 -667 926
rect -663 893 -659 900
rect -646 893 -643 935
rect -692 889 -670 893
rect -663 889 -643 893
rect -636 893 -632 944
rect -621 926 -607 930
rect -620 920 -616 926
rect -612 893 -608 900
rect -595 897 -591 940
rect -584 936 -581 948
rect -547 944 -543 962
rect -513 952 -510 958
rect -519 948 -510 952
rect -555 940 -543 944
rect -547 936 -543 940
rect -584 932 -575 936
rect -547 932 -539 936
rect -584 929 -581 932
rect -513 930 -510 948
rect -478 954 -475 966
rect -441 962 -437 976
rect -413 966 -411 970
rect -449 958 -437 962
rect -441 954 -437 958
rect -485 947 -482 954
rect -478 950 -469 954
rect -441 950 -433 954
rect -478 944 -475 950
rect -403 939 -399 976
rect -485 935 -399 939
rect -547 915 -501 919
rect -584 905 -581 908
rect -584 901 -575 905
rect -636 889 -619 893
rect -612 889 -591 893
rect -584 889 -581 901
rect -547 897 -543 915
rect -513 905 -510 907
rect -519 901 -510 905
rect -555 893 -543 897
rect -547 889 -543 893
rect -663 886 -659 889
rect -612 886 -608 889
rect -1330 871 -722 874
rect -584 885 -575 889
rect -547 885 -539 889
rect -584 879 -581 885
rect -671 870 -667 876
rect -620 870 -616 876
rect -513 870 -510 901
rect -505 893 -501 915
rect -485 901 -481 935
rect -478 905 -475 911
rect -478 901 -469 905
rect -505 889 -485 893
rect -478 889 -475 901
rect -441 897 -437 927
rect -393 905 -390 966
rect -309 948 -305 976
rect -257 952 -254 981
rect -151 970 -148 981
rect -114 976 -14 980
rect -151 966 -142 970
rect -220 962 -158 966
rect -257 948 -248 952
rect -309 944 -264 948
rect -349 926 -325 930
rect -413 901 -390 905
rect -449 893 -437 897
rect -441 889 -437 893
rect -478 885 -469 889
rect -441 885 -433 889
rect -478 879 -475 885
rect -393 870 -390 901
rect -343 920 -339 926
rect -335 893 -331 900
rect -319 893 -314 935
rect -354 889 -342 893
rect -335 889 -314 893
rect -309 893 -305 944
rect -294 926 -280 930
rect -293 920 -289 926
rect -285 893 -281 900
rect -268 897 -264 940
rect -257 936 -254 948
rect -220 944 -216 962
rect -186 952 -183 958
rect -192 948 -183 952
rect -228 940 -216 944
rect -220 936 -216 940
rect -257 932 -248 936
rect -220 932 -212 936
rect -257 929 -254 932
rect -186 930 -183 948
rect -151 954 -148 966
rect -114 962 -110 976
rect -86 966 -84 970
rect -122 958 -110 962
rect -114 954 -110 958
rect -158 947 -155 954
rect -151 950 -142 954
rect -114 950 -106 954
rect -151 944 -148 950
rect -76 939 -72 976
rect -158 935 -72 939
rect -220 915 -174 919
rect -257 905 -254 908
rect -257 901 -248 905
rect -309 889 -292 893
rect -285 889 -264 893
rect -257 889 -254 901
rect -220 897 -216 915
rect -186 905 -183 907
rect -192 901 -183 905
rect -228 893 -216 897
rect -220 889 -216 893
rect -335 886 -331 889
rect -285 886 -281 889
rect -257 885 -248 889
rect -220 885 -212 889
rect -257 879 -254 885
rect -343 870 -339 876
rect -293 870 -289 876
rect -186 870 -183 901
rect -178 893 -174 915
rect -158 901 -154 935
rect -151 905 -148 911
rect -151 901 -142 905
rect -178 889 -158 893
rect -151 889 -148 901
rect -114 897 -110 927
rect -66 905 -63 966
rect -86 901 -63 905
rect -122 893 -110 897
rect -114 889 -110 893
rect -151 885 -142 889
rect -114 885 -106 889
rect -151 879 -148 885
rect -66 870 -63 901
rect -18 898 -14 976
rect -8 906 -4 996
rect 1 982 6 1140
rect 293 1046 506 1050
rect 444 1035 487 1039
rect 407 1028 416 1032
rect 305 1024 400 1028
rect 305 994 309 1024
rect 396 1005 400 1020
rect 407 1016 410 1028
rect 444 1024 448 1035
rect 472 1028 475 1032
rect 436 1020 448 1024
rect 444 1016 448 1020
rect 353 1001 400 1005
rect 316 994 325 998
rect 273 990 309 994
rect 273 982 278 990
rect 1 977 278 982
rect 42 958 255 962
rect 193 947 236 951
rect 156 940 165 944
rect 54 936 149 940
rect 54 906 58 936
rect 145 917 149 932
rect 156 928 159 940
rect 193 936 197 947
rect 221 940 224 944
rect 185 932 197 936
rect 193 928 197 932
rect 102 913 149 917
rect 65 906 74 910
rect -8 902 58 906
rect -18 894 14 898
rect -671 867 -63 870
rect 31 826 35 902
rect 47 894 58 898
rect 65 894 68 906
rect 102 902 106 913
rect 130 906 134 910
rect 94 898 106 902
rect 102 894 106 898
rect 54 876 58 894
rect 65 890 74 894
rect 102 890 110 894
rect 145 880 149 913
rect 156 924 165 928
rect 193 924 201 928
rect 156 915 160 924
rect 156 911 205 915
rect 156 888 160 911
rect 232 906 236 947
rect 251 915 255 958
rect 274 942 278 977
rect 290 982 309 986
rect 316 982 319 994
rect 353 990 357 1001
rect 381 994 385 998
rect 345 986 357 990
rect 353 982 357 986
rect 290 968 294 982
rect 305 964 309 982
rect 316 978 325 982
rect 353 978 361 982
rect 396 968 400 1001
rect 407 1012 416 1016
rect 444 1012 452 1016
rect 407 1003 411 1012
rect 407 999 456 1003
rect 407 976 411 999
rect 483 994 487 1035
rect 502 1003 506 1046
rect 540 1002 617 1006
rect 503 994 512 998
rect 483 990 496 994
rect 483 983 496 986
rect 444 982 496 983
rect 503 982 506 994
rect 540 990 544 1002
rect 568 994 572 998
rect 532 986 544 990
rect 540 982 544 986
rect 444 979 487 982
rect 407 972 416 976
rect 305 960 400 964
rect 407 960 410 972
rect 444 968 448 979
rect 503 978 512 982
rect 540 978 548 982
rect 472 972 482 976
rect 436 964 448 968
rect 444 960 448 964
rect 407 956 416 960
rect 444 956 452 960
rect 478 953 482 972
rect 572 953 576 994
rect 293 949 576 953
rect 274 938 348 942
rect 335 918 339 920
rect 289 914 339 918
rect 252 906 261 910
rect 232 902 245 906
rect 232 895 245 898
rect 193 894 245 895
rect 252 894 255 906
rect 289 902 293 914
rect 317 906 321 910
rect 281 898 293 902
rect 289 894 293 898
rect 193 891 236 894
rect 156 884 165 888
rect 54 872 149 876
rect 156 872 159 884
rect 193 880 197 891
rect 252 890 261 894
rect 289 890 297 894
rect 221 884 231 888
rect 185 876 197 880
rect 193 872 197 876
rect 156 868 165 872
rect 193 868 201 872
rect 227 865 231 884
rect 321 865 325 906
rect 335 879 339 914
rect 344 897 348 938
rect 351 915 445 918
rect 469 915 587 918
rect 344 887 348 892
rect 362 891 365 915
rect 441 912 445 915
rect 394 894 434 898
rect 394 891 398 894
rect 362 887 368 891
rect 394 887 401 891
rect 344 883 355 887
rect 335 875 355 879
rect 362 875 365 887
rect 394 883 398 887
rect 430 883 434 894
rect 449 883 453 892
rect 456 883 473 886
rect 388 879 398 883
rect 430 879 442 883
rect 449 882 473 883
rect 449 879 459 882
rect 449 876 453 879
rect 335 871 339 875
rect 362 871 368 875
rect 421 871 427 875
rect 42 861 325 865
rect 424 863 427 871
rect 469 874 473 878
rect 480 874 483 915
rect 569 912 573 915
rect 532 893 560 896
rect 532 890 535 893
rect 526 886 535 890
rect 548 886 554 890
rect 532 882 535 886
rect 532 878 538 882
rect 551 874 554 886
rect 557 883 560 893
rect 577 883 581 892
rect 557 879 570 883
rect 577 879 592 883
rect 577 876 581 879
rect 458 870 473 874
rect 480 870 486 874
rect 548 870 554 874
rect 441 863 445 866
rect 351 860 445 863
rect 42 854 136 857
rect 53 830 56 854
rect 132 851 136 854
rect 85 833 125 837
rect 85 830 89 833
rect 53 826 59 830
rect 85 826 92 830
rect 31 822 46 826
rect 23 814 46 818
rect 53 814 56 826
rect 85 822 89 826
rect 121 822 125 833
rect 140 822 144 831
rect 153 846 446 850
rect 458 850 462 870
rect 551 863 554 870
rect 569 863 573 866
rect 469 860 581 863
rect 451 846 462 850
rect 153 822 157 846
rect 588 833 592 879
rect 274 829 368 832
rect 79 818 89 822
rect 121 818 133 822
rect 140 818 264 822
rect 140 815 144 818
rect 53 810 59 814
rect 112 810 118 814
rect 115 802 118 810
rect 132 802 136 805
rect 42 799 136 802
rect 260 801 264 818
rect 285 805 288 829
rect 364 826 368 829
rect 544 829 592 833
rect 317 808 357 812
rect 317 805 321 808
rect 285 801 291 805
rect 317 801 324 805
rect 260 797 278 801
rect 264 789 278 793
rect 285 789 288 801
rect 317 797 321 801
rect 353 797 357 808
rect 398 822 535 825
rect 372 797 376 806
rect 383 800 402 804
rect 383 797 387 800
rect 311 793 321 797
rect 353 793 365 797
rect 372 793 387 797
rect 372 790 376 793
rect 390 792 402 796
rect 390 790 394 792
rect 41 778 254 782
rect -703 767 13 771
rect -1186 752 -912 755
rect -1186 749 -1183 752
rect -916 749 -912 752
rect -1336 746 -1134 749
rect -1243 717 -1240 746
rect -1137 735 -1134 746
rect -916 746 -807 749
rect -1100 741 -964 745
rect -1137 731 -1128 735
rect -1206 727 -1144 731
rect -1243 713 -1234 717
rect -1351 709 -1250 713
rect -1336 691 -1316 695
rect -1330 685 -1326 691
rect -1322 658 -1318 665
rect -1305 658 -1302 700
rect -1351 654 -1329 658
rect -1322 654 -1302 658
rect -1295 658 -1291 709
rect -1280 691 -1266 695
rect -1279 685 -1275 691
rect -1271 658 -1267 665
rect -1254 662 -1250 705
rect -1243 701 -1240 713
rect -1206 709 -1202 727
rect -1172 717 -1169 723
rect -1178 713 -1169 717
rect -1214 705 -1202 709
rect -1206 701 -1202 705
rect -1243 697 -1234 701
rect -1206 697 -1198 701
rect -1243 694 -1240 697
rect -1172 695 -1169 713
rect -1137 719 -1134 731
rect -1100 727 -1096 741
rect -1072 731 -1070 735
rect -1108 723 -1096 727
rect -1100 719 -1096 723
rect -1144 712 -1141 719
rect -1137 715 -1128 719
rect -1100 715 -1092 719
rect -1137 709 -1134 715
rect -1062 704 -1058 741
rect -1144 700 -1058 704
rect -1206 680 -1160 684
rect -1243 670 -1240 673
rect -1243 666 -1234 670
rect -1295 654 -1278 658
rect -1271 654 -1250 658
rect -1243 654 -1240 666
rect -1206 662 -1202 680
rect -1172 670 -1169 672
rect -1178 666 -1169 670
rect -1214 658 -1202 662
rect -1206 654 -1202 658
rect -1322 651 -1318 654
rect -1271 651 -1267 654
rect -1243 650 -1234 654
rect -1206 650 -1198 654
rect -1243 644 -1240 650
rect -1330 635 -1326 641
rect -1279 635 -1275 641
rect -1172 635 -1169 666
rect -1164 658 -1160 680
rect -1144 666 -1140 700
rect -1137 670 -1134 676
rect -1137 666 -1128 670
rect -1164 654 -1144 658
rect -1137 654 -1134 666
rect -1100 662 -1096 692
rect -1052 670 -1049 731
rect -968 713 -964 741
rect -916 717 -913 746
rect -810 735 -807 746
rect -703 745 -699 767
rect -527 751 -253 754
rect -527 748 -524 751
rect -257 748 -253 751
rect -677 745 -475 748
rect -773 741 -699 745
rect -810 731 -801 735
rect -879 727 -817 731
rect -916 713 -907 717
rect -968 709 -923 713
rect -1008 691 -984 695
rect -1072 666 -1049 670
rect -1108 658 -1096 662
rect -1100 654 -1096 658
rect -1137 650 -1128 654
rect -1100 650 -1092 654
rect -1137 644 -1134 650
rect -1052 635 -1049 666
rect -1002 685 -998 691
rect -994 658 -990 665
rect -978 658 -973 700
rect -1013 654 -1001 658
rect -994 654 -973 658
rect -968 658 -964 709
rect -953 691 -939 695
rect -952 685 -948 691
rect -944 658 -940 665
rect -927 662 -923 705
rect -916 701 -913 713
rect -879 709 -875 727
rect -845 717 -842 723
rect -851 713 -842 717
rect -887 705 -875 709
rect -879 701 -875 705
rect -916 697 -907 701
rect -879 697 -871 701
rect -916 694 -913 697
rect -845 695 -842 713
rect -810 719 -807 731
rect -773 727 -769 741
rect -745 731 -743 735
rect -781 723 -769 727
rect -773 719 -769 723
rect -817 712 -814 719
rect -810 715 -801 719
rect -773 715 -765 719
rect -810 709 -807 715
rect -735 704 -731 741
rect -817 700 -731 704
rect -879 680 -833 684
rect -916 670 -913 673
rect -916 666 -907 670
rect -968 654 -951 658
rect -944 654 -923 658
rect -916 654 -913 666
rect -879 662 -875 680
rect -845 670 -842 672
rect -851 666 -842 670
rect -887 658 -875 662
rect -879 654 -875 658
rect -994 651 -990 654
rect -944 651 -940 654
rect -916 650 -907 654
rect -879 650 -871 654
rect -916 644 -913 650
rect -1002 635 -998 641
rect -952 635 -948 641
rect -845 635 -842 666
rect -837 658 -833 680
rect -817 666 -813 700
rect -810 670 -807 676
rect -810 666 -801 670
rect -837 654 -817 658
rect -810 654 -807 666
rect -773 662 -769 692
rect -725 670 -722 731
rect -584 716 -581 745
rect -478 734 -475 745
rect -257 745 -148 748
rect -441 740 -305 744
rect -478 730 -469 734
rect -547 726 -485 730
rect -584 712 -575 716
rect -692 708 -591 712
rect -677 690 -657 694
rect -745 666 -722 670
rect -781 658 -769 662
rect -773 654 -769 658
rect -810 650 -801 654
rect -773 650 -765 654
rect -810 644 -807 650
rect -725 635 -722 666
rect -671 684 -667 690
rect -663 657 -659 664
rect -646 657 -643 699
rect -692 653 -670 657
rect -663 653 -643 657
rect -636 657 -632 708
rect -621 690 -607 694
rect -620 684 -616 690
rect -612 657 -608 664
rect -595 661 -591 704
rect -584 700 -581 712
rect -547 708 -543 726
rect -513 716 -510 722
rect -519 712 -510 716
rect -555 704 -543 708
rect -547 700 -543 704
rect -584 696 -575 700
rect -547 696 -539 700
rect -584 693 -581 696
rect -513 694 -510 712
rect -478 718 -475 730
rect -441 726 -437 740
rect -413 730 -411 734
rect -449 722 -437 726
rect -441 718 -437 722
rect -485 711 -482 718
rect -478 714 -469 718
rect -441 714 -433 718
rect -478 708 -475 714
rect -403 703 -399 740
rect -485 699 -399 703
rect -547 679 -501 683
rect -584 669 -581 672
rect -584 665 -575 669
rect -636 653 -619 657
rect -612 653 -591 657
rect -584 653 -581 665
rect -547 661 -543 679
rect -513 669 -510 671
rect -519 665 -510 669
rect -555 657 -543 661
rect -547 653 -543 657
rect -663 650 -659 653
rect -612 650 -608 653
rect -1330 632 -722 635
rect -584 649 -575 653
rect -547 649 -539 653
rect -584 643 -581 649
rect -671 634 -667 640
rect -620 634 -616 640
rect -513 634 -510 665
rect -505 657 -501 679
rect -485 665 -481 699
rect -478 669 -475 675
rect -478 665 -469 669
rect -505 653 -485 657
rect -478 653 -475 665
rect -441 661 -437 691
rect -393 669 -390 730
rect -309 712 -305 740
rect -257 716 -254 745
rect -151 734 -148 745
rect -114 740 -40 744
rect -151 730 -142 734
rect -220 726 -158 730
rect -257 712 -248 716
rect -309 708 -264 712
rect -349 690 -325 694
rect -413 665 -390 669
rect -449 657 -437 661
rect -441 653 -437 657
rect -478 649 -469 653
rect -441 649 -433 653
rect -478 643 -475 649
rect -393 634 -390 665
rect -343 684 -339 690
rect -335 657 -331 664
rect -319 657 -314 699
rect -354 653 -342 657
rect -335 653 -314 657
rect -309 657 -305 708
rect -294 690 -280 694
rect -293 684 -289 690
rect -285 657 -281 664
rect -268 661 -264 704
rect -257 700 -254 712
rect -220 708 -216 726
rect -186 716 -183 722
rect -192 712 -183 716
rect -228 704 -216 708
rect -220 700 -216 704
rect -257 696 -248 700
rect -220 696 -212 700
rect -257 693 -254 696
rect -186 694 -183 712
rect -151 718 -148 730
rect -114 726 -110 740
rect -86 730 -84 734
rect -122 722 -110 726
rect -114 718 -110 722
rect -158 711 -155 718
rect -151 714 -142 718
rect -114 714 -106 718
rect -151 708 -148 714
rect -76 703 -72 740
rect -158 699 -72 703
rect -220 679 -174 683
rect -257 669 -254 672
rect -257 665 -248 669
rect -309 653 -292 657
rect -285 653 -264 657
rect -257 653 -254 665
rect -220 661 -216 679
rect -186 669 -183 671
rect -192 665 -183 669
rect -228 657 -216 661
rect -220 653 -216 657
rect -335 650 -331 653
rect -285 650 -281 653
rect -257 649 -248 653
rect -220 649 -212 653
rect -257 643 -254 649
rect -343 634 -339 640
rect -293 634 -289 640
rect -186 634 -183 665
rect -178 657 -174 679
rect -158 665 -154 699
rect -151 669 -148 675
rect -151 665 -142 669
rect -178 653 -158 657
rect -151 653 -148 665
rect -114 661 -110 691
rect -66 669 -63 730
rect -44 718 -40 740
rect 9 726 13 767
rect 192 767 235 771
rect 155 760 164 764
rect 53 756 148 760
rect 53 726 57 756
rect 144 737 148 752
rect 155 748 158 760
rect 192 756 196 767
rect 220 760 223 764
rect 184 752 196 756
rect 192 748 196 752
rect 101 733 148 737
rect 64 726 73 730
rect 9 722 57 726
rect -44 714 13 718
rect -86 665 -63 669
rect -122 657 -110 661
rect -114 653 -110 657
rect -151 649 -142 653
rect -114 649 -106 653
rect -151 643 -148 649
rect -66 634 -63 665
rect 30 646 34 722
rect 46 714 57 718
rect 64 714 67 726
rect 101 722 105 733
rect 129 726 133 730
rect 93 718 105 722
rect 101 714 105 718
rect 53 696 57 714
rect 64 710 73 714
rect 101 710 109 714
rect 144 700 148 733
rect 155 744 164 748
rect 192 744 200 748
rect 155 735 159 744
rect 155 731 204 735
rect 155 708 159 731
rect 231 726 235 767
rect 250 735 254 778
rect 264 764 268 789
rect 285 785 291 789
rect 344 785 350 789
rect 347 777 350 785
rect 384 786 394 790
rect 364 777 368 780
rect 274 774 368 777
rect 264 760 338 764
rect 334 738 338 760
rect 384 747 388 786
rect 398 757 402 788
rect 409 784 412 822
rect 517 819 521 822
rect 481 811 511 814
rect 481 808 484 811
rect 475 804 487 808
rect 481 792 484 804
rect 500 800 503 808
rect 497 796 503 800
rect 481 788 487 792
rect 500 784 503 796
rect 508 790 511 811
rect 525 790 529 799
rect 508 786 518 790
rect 525 786 533 790
rect 409 780 415 784
rect 497 780 503 784
rect 525 783 529 786
rect 409 774 412 780
rect 500 770 503 780
rect 517 770 521 773
rect 426 767 529 770
rect 398 753 493 757
rect 384 743 481 747
rect 288 734 343 738
rect 357 736 474 739
rect 251 726 260 730
rect 231 722 244 726
rect 231 715 244 718
rect 192 714 244 715
rect 251 714 254 726
rect 288 722 292 734
rect 316 726 320 730
rect 280 718 292 722
rect 288 714 292 718
rect 192 711 235 714
rect 155 704 164 708
rect 53 692 148 696
rect 155 692 158 704
rect 192 700 196 711
rect 251 710 260 714
rect 288 710 296 714
rect 220 704 230 708
rect 184 696 196 700
rect 192 692 196 696
rect 155 688 164 692
rect 192 688 200 692
rect 226 685 230 704
rect 288 697 292 710
rect 320 685 324 726
rect 339 719 343 734
rect 339 715 361 719
rect 368 715 371 736
rect 456 733 460 736
rect 400 726 450 729
rect 400 723 403 726
rect 394 719 406 723
rect 331 711 335 712
rect 368 711 374 715
rect 331 707 361 711
rect 349 699 361 703
rect 368 699 371 711
rect 399 707 403 719
rect 394 703 403 707
rect 447 704 450 726
rect 464 704 468 713
rect 477 704 481 743
rect 447 700 457 704
rect 464 700 481 704
rect 368 695 374 699
rect 436 695 442 699
rect 464 697 468 700
rect 41 681 324 685
rect 439 684 442 695
rect 456 684 460 687
rect 357 681 468 684
rect 41 674 135 677
rect 52 650 55 674
rect 131 671 135 674
rect 489 672 493 753
rect 544 751 548 829
rect 84 653 124 657
rect 84 650 88 653
rect 52 646 58 650
rect 84 646 91 650
rect 30 642 45 646
rect 22 634 45 638
rect 52 634 55 646
rect 84 642 88 646
rect 120 642 124 653
rect 139 642 143 651
rect 152 668 493 672
rect 152 642 156 668
rect 173 651 386 655
rect 78 638 88 642
rect 120 638 132 642
rect 139 638 156 642
rect 324 640 367 644
rect 139 635 143 638
rect -671 631 -63 634
rect 52 630 58 634
rect 111 630 117 634
rect 114 622 117 630
rect 287 633 296 637
rect 185 629 280 633
rect 131 622 135 625
rect 41 619 135 622
rect 185 599 189 629
rect 276 610 280 625
rect 287 621 290 633
rect 324 629 328 640
rect 352 633 355 637
rect 316 625 328 629
rect 324 621 328 625
rect 233 606 280 610
rect 196 599 205 603
rect 167 595 189 599
rect 167 587 189 591
rect 196 587 199 599
rect 233 595 237 606
rect 261 599 265 603
rect 225 591 237 595
rect 233 587 237 591
rect -703 546 15 550
rect -1186 538 -912 541
rect -1186 535 -1183 538
rect -916 535 -912 538
rect -1336 532 -1134 535
rect -1243 503 -1240 532
rect -1137 521 -1134 532
rect -916 532 -807 535
rect -1100 527 -964 531
rect -1137 517 -1128 521
rect -1206 513 -1144 517
rect -1243 499 -1234 503
rect -1351 495 -1250 499
rect -1336 477 -1316 481
rect -1330 471 -1326 477
rect -1322 444 -1318 451
rect -1305 444 -1302 486
rect -1351 440 -1329 444
rect -1322 440 -1302 444
rect -1295 444 -1291 495
rect -1280 477 -1266 481
rect -1279 471 -1275 477
rect -1271 444 -1267 451
rect -1254 448 -1250 491
rect -1243 487 -1240 499
rect -1206 495 -1202 513
rect -1172 503 -1169 509
rect -1178 499 -1169 503
rect -1214 491 -1202 495
rect -1206 487 -1202 491
rect -1243 483 -1234 487
rect -1206 483 -1198 487
rect -1243 480 -1240 483
rect -1172 481 -1169 499
rect -1137 505 -1134 517
rect -1100 513 -1096 527
rect -1072 517 -1070 521
rect -1108 509 -1096 513
rect -1100 505 -1096 509
rect -1144 498 -1141 505
rect -1137 501 -1128 505
rect -1100 501 -1092 505
rect -1137 495 -1134 501
rect -1062 490 -1058 527
rect -1144 486 -1058 490
rect -1206 466 -1160 470
rect -1243 456 -1240 459
rect -1243 452 -1234 456
rect -1295 440 -1278 444
rect -1271 440 -1250 444
rect -1243 440 -1240 452
rect -1206 448 -1202 466
rect -1172 456 -1169 458
rect -1178 452 -1169 456
rect -1214 444 -1202 448
rect -1206 440 -1202 444
rect -1322 437 -1318 440
rect -1271 437 -1267 440
rect -1243 436 -1234 440
rect -1206 436 -1198 440
rect -1243 430 -1240 436
rect -1330 421 -1326 427
rect -1279 421 -1275 427
rect -1172 421 -1169 452
rect -1164 444 -1160 466
rect -1144 452 -1140 486
rect -1137 456 -1134 462
rect -1137 452 -1128 456
rect -1164 440 -1144 444
rect -1137 440 -1134 452
rect -1100 448 -1096 478
rect -1052 456 -1049 517
rect -968 499 -964 527
rect -916 503 -913 532
rect -810 521 -807 532
rect -703 531 -699 546
rect -527 537 -253 540
rect -527 534 -524 537
rect -257 534 -253 537
rect -677 531 -475 534
rect -773 527 -699 531
rect -810 517 -801 521
rect -879 513 -817 517
rect -916 499 -907 503
rect -968 495 -923 499
rect -1008 477 -984 481
rect -1072 452 -1049 456
rect -1108 444 -1096 448
rect -1100 440 -1096 444
rect -1137 436 -1128 440
rect -1100 436 -1092 440
rect -1137 430 -1134 436
rect -1052 421 -1049 452
rect -1002 471 -998 477
rect -994 444 -990 451
rect -978 444 -973 486
rect -1013 440 -1001 444
rect -994 440 -973 444
rect -968 444 -964 495
rect -953 477 -939 481
rect -952 471 -948 477
rect -944 444 -940 451
rect -927 448 -923 491
rect -916 487 -913 499
rect -879 495 -875 513
rect -845 503 -842 509
rect -851 499 -842 503
rect -887 491 -875 495
rect -879 487 -875 491
rect -916 483 -907 487
rect -879 483 -871 487
rect -916 480 -913 483
rect -845 481 -842 499
rect -810 505 -807 517
rect -773 513 -769 527
rect -745 517 -743 521
rect -781 509 -769 513
rect -773 505 -769 509
rect -817 498 -814 505
rect -810 501 -801 505
rect -773 501 -765 505
rect -810 495 -807 501
rect -735 490 -731 527
rect -817 486 -731 490
rect -879 466 -833 470
rect -916 456 -913 459
rect -916 452 -907 456
rect -968 440 -951 444
rect -944 440 -923 444
rect -916 440 -913 452
rect -879 448 -875 466
rect -845 456 -842 458
rect -851 452 -842 456
rect -887 444 -875 448
rect -879 440 -875 444
rect -994 437 -990 440
rect -944 437 -940 440
rect -916 436 -907 440
rect -879 436 -871 440
rect -916 430 -913 436
rect -1002 421 -998 427
rect -952 421 -948 427
rect -845 421 -842 452
rect -837 444 -833 466
rect -817 452 -813 486
rect -810 456 -807 462
rect -810 452 -801 456
rect -837 440 -817 444
rect -810 440 -807 452
rect -773 448 -769 478
rect -725 456 -722 517
rect -584 502 -581 531
rect -478 520 -475 531
rect -257 531 -148 534
rect -441 526 -305 530
rect -478 516 -469 520
rect -547 512 -485 516
rect -584 498 -575 502
rect -692 494 -591 498
rect -677 476 -657 480
rect -745 452 -722 456
rect -781 444 -769 448
rect -773 440 -769 444
rect -810 436 -801 440
rect -773 436 -765 440
rect -810 430 -807 436
rect -725 421 -722 452
rect -671 470 -667 476
rect -663 443 -659 450
rect -646 443 -643 485
rect -692 439 -670 443
rect -663 439 -643 443
rect -636 443 -632 494
rect -621 476 -607 480
rect -620 470 -616 476
rect -612 443 -608 450
rect -595 447 -591 490
rect -584 486 -581 498
rect -547 494 -543 512
rect -513 502 -510 508
rect -519 498 -510 502
rect -555 490 -543 494
rect -547 486 -543 490
rect -584 482 -575 486
rect -547 482 -539 486
rect -584 479 -581 482
rect -513 480 -510 498
rect -478 504 -475 516
rect -441 512 -437 526
rect -413 516 -411 520
rect -449 508 -437 512
rect -441 504 -437 508
rect -485 497 -482 504
rect -478 500 -469 504
rect -441 500 -433 504
rect -478 494 -475 500
rect -403 489 -399 526
rect -485 485 -399 489
rect -547 465 -501 469
rect -584 455 -581 458
rect -584 451 -575 455
rect -636 439 -619 443
rect -612 439 -591 443
rect -584 439 -581 451
rect -547 447 -543 465
rect -513 455 -510 457
rect -519 451 -510 455
rect -555 443 -543 447
rect -547 439 -543 443
rect -663 436 -659 439
rect -612 436 -608 439
rect -1330 418 -722 421
rect -584 435 -575 439
rect -547 435 -539 439
rect -584 429 -581 435
rect -671 420 -667 426
rect -620 420 -616 426
rect -513 420 -510 451
rect -505 443 -501 465
rect -485 451 -481 485
rect -478 455 -475 461
rect -478 451 -469 455
rect -505 439 -485 443
rect -478 439 -475 451
rect -441 447 -437 477
rect -393 455 -390 516
rect -309 498 -305 526
rect -257 502 -254 531
rect -151 520 -148 531
rect -114 526 -40 530
rect -151 516 -142 520
rect -220 512 -158 516
rect -257 498 -248 502
rect -309 494 -264 498
rect -349 476 -325 480
rect -413 451 -390 455
rect -449 443 -437 447
rect -441 439 -437 443
rect -478 435 -469 439
rect -441 435 -433 439
rect -478 429 -475 435
rect -393 420 -390 451
rect -343 470 -339 476
rect -335 443 -331 450
rect -319 443 -314 485
rect -354 439 -342 443
rect -335 439 -314 443
rect -309 443 -305 494
rect -294 476 -280 480
rect -293 470 -289 476
rect -285 443 -281 450
rect -268 447 -264 490
rect -257 486 -254 498
rect -220 494 -216 512
rect -186 502 -183 508
rect -192 498 -183 502
rect -228 490 -216 494
rect -220 486 -216 490
rect -257 482 -248 486
rect -220 482 -212 486
rect -257 479 -254 482
rect -186 480 -183 498
rect -151 504 -148 516
rect -114 512 -110 526
rect -86 516 -84 520
rect -122 508 -110 512
rect -114 504 -110 508
rect -158 497 -155 504
rect -151 500 -142 504
rect -114 500 -106 504
rect -151 494 -148 500
rect -76 489 -72 526
rect -158 485 -72 489
rect -220 465 -174 469
rect -257 455 -254 458
rect -257 451 -248 455
rect -309 439 -292 443
rect -285 439 -264 443
rect -257 439 -254 451
rect -220 447 -216 465
rect -186 455 -183 457
rect -192 451 -183 455
rect -228 443 -216 447
rect -220 439 -216 443
rect -335 436 -331 439
rect -285 436 -281 439
rect -257 435 -248 439
rect -220 435 -212 439
rect -257 429 -254 435
rect -343 420 -339 426
rect -293 420 -289 426
rect -186 420 -183 451
rect -178 443 -174 465
rect -158 451 -154 485
rect -151 455 -148 461
rect -151 451 -142 455
rect -178 439 -158 443
rect -151 439 -148 451
rect -114 447 -110 477
rect -66 455 -63 516
rect -44 464 -40 526
rect 11 472 15 546
rect 167 544 170 587
rect 185 569 189 587
rect 196 583 205 587
rect 233 583 241 587
rect 276 573 280 606
rect 287 617 296 621
rect 324 617 332 621
rect 287 608 291 617
rect 287 604 336 608
rect 287 581 291 604
rect 363 599 367 640
rect 382 608 386 651
rect 420 607 474 611
rect 383 599 392 603
rect 363 595 376 599
rect 363 588 376 591
rect 324 587 376 588
rect 383 587 386 599
rect 420 595 424 607
rect 448 599 452 603
rect 412 591 424 595
rect 420 587 424 591
rect 324 584 367 587
rect 287 577 296 581
rect 185 565 280 569
rect 287 565 290 577
rect 324 573 328 584
rect 383 583 392 587
rect 420 583 428 587
rect 352 577 362 581
rect 316 569 328 573
rect 324 565 328 569
rect 287 561 296 565
rect 324 561 332 565
rect 358 558 362 577
rect 452 558 456 599
rect 173 554 456 558
rect 470 557 474 607
rect 489 564 493 668
rect 502 747 548 751
rect 502 544 506 747
rect 613 731 617 1002
rect 635 895 638 1162
rect 717 1162 746 1165
rect 677 1114 681 1155
rect 685 1151 728 1155
rect 695 1130 699 1139
rect 732 1138 736 1155
rect 725 1134 739 1138
rect 695 1126 705 1130
rect 755 1130 758 1233
rect 783 1268 823 1271
rect 783 1166 786 1268
rect 828 1265 832 1343
rect 862 1333 866 1353
rect 878 1309 882 1313
rect 840 1305 882 1309
rect 870 1297 874 1305
rect 862 1271 866 1277
rect 878 1271 882 1277
rect 856 1268 888 1271
rect 813 1261 820 1264
rect 801 1203 805 1261
rect 828 1261 866 1265
rect 874 1245 878 1261
rect 848 1241 878 1245
rect 809 1233 837 1236
rect 815 1227 819 1233
rect 831 1203 835 1207
rect 801 1199 835 1203
rect 848 1203 852 1241
rect 897 1236 900 1353
rect 927 1347 931 1379
rect 941 1353 1040 1356
rect 927 1343 972 1347
rect 927 1309 931 1343
rect 937 1333 941 1335
rect 953 1309 957 1313
rect 927 1305 957 1309
rect 945 1297 949 1305
rect 937 1271 941 1277
rect 953 1271 957 1277
rect 860 1233 900 1236
rect 862 1227 866 1233
rect 878 1203 882 1207
rect 848 1199 882 1203
rect 823 1191 827 1199
rect 870 1191 874 1199
rect 695 1125 699 1126
rect 732 1114 736 1127
rect 749 1126 758 1130
rect 645 1110 736 1114
rect 645 1020 649 1110
rect 690 1100 736 1105
rect 695 1080 699 1094
rect 732 1088 736 1100
rect 725 1084 739 1088
rect 695 1076 705 1080
rect 755 1080 758 1126
rect 695 1070 699 1076
rect 732 1065 736 1077
rect 749 1076 758 1080
rect 755 1029 758 1076
rect 659 1026 758 1029
rect 645 1016 690 1020
rect 645 982 649 1016
rect 655 1006 659 1008
rect 671 982 675 986
rect 645 978 675 982
rect 663 970 667 978
rect 655 944 659 950
rect 671 944 675 950
rect 641 941 681 944
rect 641 895 644 941
rect 686 938 690 1016
rect 720 1006 724 1026
rect 736 982 740 986
rect 698 978 740 982
rect 728 970 732 978
rect 720 944 724 950
rect 736 944 740 950
rect 714 941 746 944
rect 671 934 678 937
rect 635 892 644 895
rect 641 838 644 892
rect 659 876 663 934
rect 686 934 724 938
rect 732 918 736 934
rect 706 914 736 918
rect 667 906 695 909
rect 673 900 677 906
rect 689 876 693 880
rect 659 872 693 876
rect 706 876 710 914
rect 755 909 758 1026
rect 718 906 758 909
rect 720 900 724 906
rect 736 876 740 880
rect 706 872 740 876
rect 681 864 685 872
rect 728 864 732 872
rect 673 838 677 844
rect 689 838 693 844
rect 720 838 724 844
rect 736 838 740 844
rect 641 835 696 838
rect 641 742 644 835
rect 717 835 746 838
rect 677 787 681 828
rect 685 824 728 828
rect 695 803 699 812
rect 732 811 736 828
rect 725 807 739 811
rect 695 799 705 803
rect 755 803 758 906
rect 777 1165 786 1166
rect 815 1165 819 1171
rect 831 1165 835 1171
rect 862 1165 866 1171
rect 878 1165 882 1171
rect 777 1162 838 1165
rect 777 895 780 1162
rect 859 1162 888 1165
rect 819 1114 823 1155
rect 827 1151 870 1155
rect 837 1130 841 1139
rect 874 1138 878 1155
rect 867 1134 881 1138
rect 837 1126 847 1130
rect 897 1130 900 1233
rect 923 1268 963 1271
rect 923 1166 926 1268
rect 968 1265 972 1343
rect 1002 1333 1006 1353
rect 1018 1309 1022 1313
rect 980 1305 1022 1309
rect 1010 1297 1014 1305
rect 1002 1271 1006 1277
rect 1018 1271 1022 1277
rect 996 1268 1028 1271
rect 953 1261 960 1264
rect 941 1203 945 1261
rect 968 1261 1006 1265
rect 1014 1245 1018 1261
rect 988 1241 1018 1245
rect 949 1233 977 1236
rect 955 1227 959 1233
rect 971 1203 975 1207
rect 941 1199 975 1203
rect 988 1203 992 1241
rect 1037 1236 1040 1353
rect 1072 1347 1076 1379
rect 1086 1353 1185 1356
rect 1072 1343 1117 1347
rect 1072 1309 1076 1343
rect 1082 1333 1086 1335
rect 1098 1309 1102 1313
rect 1072 1305 1102 1309
rect 1090 1297 1094 1305
rect 1082 1271 1086 1277
rect 1098 1271 1102 1277
rect 1000 1233 1040 1236
rect 1002 1227 1006 1233
rect 1018 1203 1022 1207
rect 988 1199 1022 1203
rect 963 1191 967 1199
rect 1010 1191 1014 1199
rect 837 1125 841 1126
rect 874 1114 878 1127
rect 891 1126 900 1130
rect 787 1110 878 1114
rect 787 1020 791 1110
rect 832 1100 878 1105
rect 837 1080 841 1094
rect 874 1088 878 1100
rect 867 1084 881 1088
rect 837 1076 847 1080
rect 897 1080 900 1126
rect 837 1070 841 1076
rect 874 1065 878 1077
rect 891 1076 900 1080
rect 897 1029 900 1076
rect 801 1026 900 1029
rect 787 1016 832 1020
rect 787 982 791 1016
rect 797 1006 801 1008
rect 813 982 817 986
rect 787 978 817 982
rect 805 970 809 978
rect 797 944 801 950
rect 813 944 817 950
rect 783 941 823 944
rect 783 895 786 941
rect 828 938 832 1016
rect 862 1006 866 1026
rect 878 982 882 986
rect 840 978 882 982
rect 870 970 874 978
rect 862 944 866 950
rect 878 944 882 950
rect 856 941 888 944
rect 813 934 820 937
rect 777 892 786 895
rect 695 798 699 799
rect 732 787 736 800
rect 749 799 758 803
rect 677 783 736 787
rect 677 731 681 783
rect 690 773 736 776
rect 695 752 699 762
rect 732 760 736 773
rect 725 756 739 760
rect 695 748 705 752
rect 755 752 758 799
rect 695 742 699 748
rect 613 727 681 731
rect 732 727 736 749
rect 749 748 758 752
rect 783 838 786 892
rect 801 876 805 934
rect 828 934 866 938
rect 874 918 878 934
rect 848 914 878 918
rect 809 906 837 909
rect 815 900 819 906
rect 831 876 835 880
rect 801 872 835 876
rect 848 876 852 914
rect 897 909 900 1026
rect 860 906 900 909
rect 862 900 866 906
rect 878 876 882 880
rect 848 872 882 876
rect 823 864 827 872
rect 870 864 874 872
rect 815 838 819 844
rect 831 838 835 844
rect 862 838 866 844
rect 878 838 882 844
rect 783 835 838 838
rect 783 742 786 835
rect 859 835 888 838
rect 819 787 823 828
rect 827 824 870 828
rect 837 803 841 812
rect 874 811 878 828
rect 867 807 881 811
rect 837 799 847 803
rect 897 803 900 906
rect 917 1165 926 1166
rect 955 1165 959 1171
rect 971 1165 975 1171
rect 1002 1165 1006 1171
rect 1018 1165 1022 1171
rect 917 1162 978 1165
rect 917 895 920 1162
rect 999 1162 1028 1165
rect 959 1114 963 1155
rect 967 1151 1010 1155
rect 977 1130 981 1139
rect 1014 1138 1018 1155
rect 1007 1134 1021 1138
rect 977 1126 987 1130
rect 1037 1130 1040 1233
rect 1068 1268 1108 1271
rect 1068 1166 1071 1268
rect 1113 1265 1117 1343
rect 1147 1333 1151 1353
rect 1163 1309 1167 1313
rect 1125 1305 1167 1309
rect 1155 1297 1159 1305
rect 1147 1271 1151 1277
rect 1163 1271 1167 1277
rect 1141 1268 1173 1271
rect 1098 1261 1105 1264
rect 1086 1203 1090 1261
rect 1113 1261 1151 1265
rect 1159 1245 1163 1261
rect 1133 1241 1163 1245
rect 1094 1233 1122 1236
rect 1100 1227 1104 1233
rect 1116 1203 1120 1207
rect 1086 1199 1120 1203
rect 1133 1203 1137 1241
rect 1182 1236 1185 1353
rect 1217 1347 1221 1379
rect 1231 1353 1330 1356
rect 1217 1343 1262 1347
rect 1217 1309 1221 1343
rect 1227 1333 1231 1335
rect 1243 1309 1247 1313
rect 1217 1305 1247 1309
rect 1235 1297 1239 1305
rect 1227 1271 1231 1277
rect 1243 1271 1247 1277
rect 1145 1233 1185 1236
rect 1147 1227 1151 1233
rect 1163 1203 1167 1207
rect 1133 1199 1167 1203
rect 1108 1191 1112 1199
rect 1155 1191 1159 1199
rect 977 1125 981 1126
rect 1014 1114 1018 1127
rect 1031 1126 1040 1130
rect 927 1110 1018 1114
rect 927 1020 931 1110
rect 972 1100 1018 1105
rect 977 1080 981 1094
rect 1014 1088 1018 1100
rect 1007 1084 1021 1088
rect 977 1076 987 1080
rect 1037 1080 1040 1126
rect 977 1070 981 1076
rect 1014 1065 1018 1077
rect 1031 1076 1040 1080
rect 1037 1029 1040 1076
rect 941 1026 1040 1029
rect 927 1016 972 1020
rect 927 982 931 1016
rect 937 1006 941 1008
rect 953 982 957 986
rect 927 978 957 982
rect 945 970 949 978
rect 937 944 941 950
rect 953 944 957 950
rect 923 941 963 944
rect 923 895 926 941
rect 968 938 972 1016
rect 1002 1006 1006 1026
rect 1018 982 1022 986
rect 980 978 1022 982
rect 1010 970 1014 978
rect 1002 944 1006 950
rect 1018 944 1022 950
rect 996 941 1028 944
rect 953 934 960 937
rect 917 892 926 895
rect 837 798 841 799
rect 874 787 878 800
rect 891 799 900 803
rect 819 783 878 787
rect 819 733 823 783
rect 832 773 878 776
rect 837 752 841 762
rect 874 760 878 773
rect 867 756 881 760
rect 837 748 847 752
rect 897 752 900 799
rect 837 742 841 748
rect 874 727 878 749
rect 891 748 900 752
rect 923 838 926 892
rect 941 876 945 934
rect 968 934 1006 938
rect 1014 918 1018 934
rect 988 914 1018 918
rect 949 906 977 909
rect 955 900 959 906
rect 971 876 975 880
rect 941 872 975 876
rect 988 876 992 914
rect 1037 909 1040 1026
rect 1000 906 1040 909
rect 1002 900 1006 906
rect 1018 876 1022 880
rect 988 872 1022 876
rect 963 864 967 872
rect 1010 864 1014 872
rect 955 838 959 844
rect 971 838 975 844
rect 1002 838 1006 844
rect 1018 838 1022 844
rect 923 835 978 838
rect 923 742 926 835
rect 999 835 1028 838
rect 959 787 963 828
rect 967 824 1010 828
rect 977 803 981 812
rect 1014 811 1018 828
rect 1007 807 1021 811
rect 977 799 987 803
rect 1037 803 1040 906
rect 1062 1165 1071 1166
rect 1100 1165 1104 1171
rect 1116 1165 1120 1171
rect 1147 1165 1151 1171
rect 1163 1165 1167 1171
rect 1062 1162 1123 1165
rect 1062 895 1065 1162
rect 1144 1162 1173 1165
rect 1104 1114 1108 1155
rect 1112 1151 1155 1155
rect 1122 1130 1126 1139
rect 1159 1138 1163 1155
rect 1152 1134 1166 1138
rect 1122 1126 1132 1130
rect 1182 1130 1185 1233
rect 1213 1268 1253 1271
rect 1213 1166 1216 1268
rect 1258 1265 1262 1343
rect 1292 1333 1296 1353
rect 1308 1309 1312 1313
rect 1270 1305 1312 1309
rect 1300 1297 1304 1305
rect 1292 1271 1296 1277
rect 1308 1271 1312 1277
rect 1286 1268 1318 1271
rect 1243 1261 1250 1264
rect 1231 1203 1235 1261
rect 1258 1261 1296 1265
rect 1304 1245 1308 1261
rect 1278 1241 1308 1245
rect 1239 1233 1267 1236
rect 1245 1227 1249 1233
rect 1261 1203 1265 1207
rect 1231 1199 1265 1203
rect 1278 1203 1282 1241
rect 1327 1236 1330 1353
rect 1362 1347 1366 1379
rect 1376 1353 1475 1356
rect 1362 1343 1407 1347
rect 1362 1309 1366 1343
rect 1372 1333 1376 1335
rect 1388 1309 1392 1313
rect 1362 1305 1392 1309
rect 1380 1297 1384 1305
rect 1372 1271 1376 1277
rect 1388 1271 1392 1277
rect 1290 1233 1330 1236
rect 1292 1227 1296 1233
rect 1308 1203 1312 1207
rect 1278 1199 1312 1203
rect 1253 1191 1257 1199
rect 1300 1191 1304 1199
rect 1122 1125 1126 1126
rect 1159 1114 1163 1127
rect 1176 1126 1185 1130
rect 1072 1110 1163 1114
rect 1072 1020 1076 1110
rect 1117 1100 1163 1105
rect 1122 1080 1126 1094
rect 1159 1088 1163 1100
rect 1152 1084 1166 1088
rect 1122 1076 1132 1080
rect 1182 1080 1185 1126
rect 1122 1070 1126 1076
rect 1159 1065 1163 1077
rect 1176 1076 1185 1080
rect 1182 1029 1185 1076
rect 1086 1026 1185 1029
rect 1072 1016 1117 1020
rect 1072 982 1076 1016
rect 1082 1006 1086 1008
rect 1098 982 1102 986
rect 1072 978 1102 982
rect 1090 970 1094 978
rect 1082 944 1086 950
rect 1098 944 1102 950
rect 1068 941 1108 944
rect 1068 895 1071 941
rect 1113 938 1117 1016
rect 1147 1006 1151 1026
rect 1163 982 1167 986
rect 1125 978 1167 982
rect 1155 970 1159 978
rect 1147 944 1151 950
rect 1163 944 1167 950
rect 1141 941 1173 944
rect 1098 934 1105 937
rect 1062 892 1071 895
rect 977 798 981 799
rect 1014 787 1018 800
rect 1031 799 1040 803
rect 959 783 1018 787
rect 532 691 745 695
rect 683 680 726 684
rect 646 673 655 677
rect 544 669 639 673
rect 544 639 548 669
rect 635 650 639 665
rect 646 661 649 673
rect 683 669 687 680
rect 711 673 714 677
rect 675 665 687 669
rect 683 661 687 665
rect 592 646 639 650
rect 555 639 564 643
rect 536 636 548 639
rect 532 635 548 636
rect 167 540 506 544
rect 518 627 548 631
rect 555 627 558 639
rect 592 635 596 646
rect 620 639 624 643
rect 584 631 596 635
rect 592 627 596 631
rect 342 532 369 535
rect 41 524 254 528
rect 192 513 235 517
rect 155 506 164 510
rect 53 502 148 506
rect 53 472 57 502
rect 144 483 148 498
rect 155 494 158 506
rect 192 502 196 513
rect 220 506 223 510
rect 184 498 196 502
rect 192 494 196 498
rect 101 479 148 483
rect 64 472 73 476
rect 11 468 57 472
rect -44 460 13 464
rect -86 451 -63 455
rect -122 443 -110 447
rect -114 439 -110 443
rect -151 435 -142 439
rect -114 435 -106 439
rect -151 429 -148 435
rect -66 420 -63 451
rect -671 417 -63 420
rect 30 392 34 468
rect 46 460 57 464
rect 64 460 67 472
rect 101 468 105 479
rect 129 472 133 476
rect 93 464 105 468
rect 101 460 105 464
rect 53 442 57 460
rect 64 456 73 460
rect 101 456 109 460
rect 144 446 148 479
rect 155 490 164 494
rect 192 490 200 494
rect 155 481 159 490
rect 155 477 204 481
rect 155 454 159 477
rect 231 472 235 513
rect 250 481 254 524
rect 342 512 345 532
rect 471 521 474 531
rect 518 527 522 627
rect 544 609 548 627
rect 555 623 564 627
rect 592 623 600 627
rect 635 613 639 646
rect 646 657 655 661
rect 683 657 691 661
rect 646 648 650 657
rect 646 644 695 648
rect 646 621 650 644
rect 722 639 726 680
rect 741 648 745 691
rect 779 650 894 651
rect 959 650 963 783
rect 972 773 1018 776
rect 977 752 981 762
rect 1014 760 1018 773
rect 1007 756 1021 760
rect 977 748 987 752
rect 1037 752 1040 799
rect 977 742 981 748
rect 1014 727 1018 749
rect 1031 748 1040 752
rect 1068 838 1071 892
rect 1086 876 1090 934
rect 1113 934 1151 938
rect 1159 918 1163 934
rect 1133 914 1163 918
rect 1094 906 1122 909
rect 1100 900 1104 906
rect 1116 876 1120 880
rect 1086 872 1120 876
rect 1133 876 1137 914
rect 1182 909 1185 1026
rect 1145 906 1185 909
rect 1147 900 1151 906
rect 1163 876 1167 880
rect 1133 872 1167 876
rect 1108 864 1112 872
rect 1155 864 1159 872
rect 1100 838 1104 844
rect 1116 838 1120 844
rect 1147 838 1151 844
rect 1163 838 1167 844
rect 1068 835 1123 838
rect 1068 742 1071 835
rect 1144 835 1173 838
rect 1104 787 1108 828
rect 1112 824 1155 828
rect 1122 803 1126 812
rect 1159 811 1163 828
rect 1152 807 1166 811
rect 1122 799 1132 803
rect 1182 803 1185 906
rect 1207 1165 1216 1166
rect 1245 1165 1249 1171
rect 1261 1165 1265 1171
rect 1292 1165 1296 1171
rect 1308 1165 1312 1171
rect 1207 1162 1268 1165
rect 1207 895 1210 1162
rect 1289 1162 1318 1165
rect 1249 1114 1253 1155
rect 1257 1151 1300 1155
rect 1267 1130 1271 1139
rect 1304 1138 1308 1155
rect 1297 1134 1311 1138
rect 1267 1126 1277 1130
rect 1327 1130 1330 1233
rect 1358 1268 1398 1271
rect 1358 1166 1361 1268
rect 1403 1265 1407 1343
rect 1437 1333 1441 1353
rect 1453 1309 1457 1313
rect 1415 1305 1457 1309
rect 1445 1297 1449 1305
rect 1437 1271 1441 1277
rect 1453 1271 1457 1277
rect 1431 1268 1463 1271
rect 1388 1261 1395 1264
rect 1376 1203 1380 1261
rect 1403 1261 1441 1265
rect 1449 1245 1453 1261
rect 1423 1241 1453 1245
rect 1384 1233 1412 1236
rect 1390 1227 1394 1233
rect 1406 1203 1410 1207
rect 1376 1199 1410 1203
rect 1423 1203 1427 1241
rect 1472 1236 1475 1353
rect 1435 1233 1475 1236
rect 1437 1227 1441 1233
rect 1453 1203 1457 1207
rect 1423 1199 1457 1203
rect 1398 1191 1402 1199
rect 1445 1191 1449 1199
rect 1267 1125 1271 1126
rect 1304 1114 1308 1127
rect 1321 1126 1330 1130
rect 1217 1110 1308 1114
rect 1217 1020 1221 1110
rect 1262 1100 1308 1105
rect 1267 1080 1271 1094
rect 1304 1088 1308 1100
rect 1297 1084 1311 1088
rect 1267 1076 1277 1080
rect 1327 1080 1330 1126
rect 1267 1070 1271 1076
rect 1304 1065 1308 1077
rect 1321 1076 1330 1080
rect 1327 1029 1330 1076
rect 1231 1026 1330 1029
rect 1217 1016 1262 1020
rect 1217 982 1221 1016
rect 1227 1006 1231 1008
rect 1243 982 1247 986
rect 1217 978 1247 982
rect 1235 970 1239 978
rect 1227 944 1231 950
rect 1243 944 1247 950
rect 1213 941 1253 944
rect 1213 895 1216 941
rect 1258 938 1262 1016
rect 1292 1006 1296 1026
rect 1308 982 1312 986
rect 1270 978 1312 982
rect 1300 970 1304 978
rect 1292 944 1296 950
rect 1308 944 1312 950
rect 1286 941 1318 944
rect 1243 934 1250 937
rect 1207 892 1216 895
rect 1122 798 1126 799
rect 1159 787 1163 800
rect 1176 799 1185 803
rect 1104 783 1163 787
rect 1104 722 1108 783
rect 1117 773 1163 776
rect 1122 752 1126 762
rect 1159 760 1163 773
rect 1152 756 1166 760
rect 1122 748 1132 752
rect 1182 752 1185 799
rect 1122 742 1126 748
rect 1159 727 1163 749
rect 1176 748 1185 752
rect 1213 838 1216 892
rect 1231 876 1235 934
rect 1258 934 1296 938
rect 1304 918 1308 934
rect 1278 914 1308 918
rect 1239 906 1267 909
rect 1245 900 1249 906
rect 1261 876 1265 880
rect 1231 872 1265 876
rect 1278 876 1282 914
rect 1327 909 1330 1026
rect 1290 906 1330 909
rect 1292 900 1296 906
rect 1308 876 1312 880
rect 1278 872 1312 876
rect 1253 864 1257 872
rect 1300 864 1304 872
rect 1245 838 1249 844
rect 1261 838 1265 844
rect 1292 838 1296 844
rect 1308 838 1312 844
rect 1213 835 1268 838
rect 1213 742 1216 835
rect 1289 835 1318 838
rect 1249 787 1253 828
rect 1257 824 1300 828
rect 1267 803 1271 812
rect 1304 811 1308 828
rect 1297 807 1311 811
rect 1267 799 1277 803
rect 1327 803 1330 906
rect 1352 1165 1361 1166
rect 1390 1165 1394 1171
rect 1406 1165 1410 1171
rect 1437 1165 1441 1171
rect 1453 1165 1457 1171
rect 1352 1162 1413 1165
rect 1352 895 1355 1162
rect 1434 1162 1463 1165
rect 1394 1114 1398 1155
rect 1402 1151 1445 1155
rect 1412 1130 1416 1139
rect 1449 1138 1453 1155
rect 1442 1134 1456 1138
rect 1412 1126 1422 1130
rect 1472 1130 1475 1233
rect 1412 1125 1416 1126
rect 1449 1114 1453 1127
rect 1466 1126 1475 1130
rect 1362 1110 1453 1114
rect 1362 1020 1366 1110
rect 1407 1100 1453 1105
rect 1412 1080 1416 1094
rect 1449 1088 1453 1100
rect 1442 1084 1456 1088
rect 1412 1076 1422 1080
rect 1472 1080 1475 1126
rect 1412 1070 1416 1076
rect 1449 1065 1453 1077
rect 1466 1076 1475 1080
rect 1472 1029 1475 1076
rect 1376 1026 1475 1029
rect 1362 1016 1407 1020
rect 1362 982 1366 1016
rect 1372 1006 1376 1008
rect 1388 982 1392 986
rect 1362 978 1392 982
rect 1380 970 1384 978
rect 1372 944 1376 950
rect 1388 944 1392 950
rect 1358 941 1398 944
rect 1358 895 1361 941
rect 1403 938 1407 1016
rect 1437 1006 1441 1026
rect 1453 982 1457 986
rect 1415 978 1457 982
rect 1445 970 1449 978
rect 1437 944 1441 950
rect 1453 944 1457 950
rect 1431 941 1463 944
rect 1388 934 1395 937
rect 1352 892 1361 895
rect 1267 798 1271 799
rect 1304 787 1308 800
rect 1321 799 1330 803
rect 1249 783 1308 787
rect 779 647 963 650
rect 742 639 751 643
rect 722 635 735 639
rect 722 628 735 631
rect 683 627 735 628
rect 742 627 745 639
rect 779 635 783 647
rect 894 646 963 647
rect 976 718 1108 722
rect 807 639 811 643
rect 976 642 980 718
rect 1249 713 1253 783
rect 1262 773 1308 776
rect 1267 752 1271 762
rect 1304 760 1308 773
rect 1297 756 1311 760
rect 1267 748 1277 752
rect 1327 752 1330 799
rect 1267 742 1271 748
rect 1304 727 1308 749
rect 1321 748 1330 752
rect 1358 838 1361 892
rect 1376 876 1380 934
rect 1403 934 1441 938
rect 1449 918 1453 934
rect 1423 914 1453 918
rect 1384 906 1412 909
rect 1390 900 1394 906
rect 1406 876 1410 880
rect 1376 872 1410 876
rect 1423 876 1427 914
rect 1472 909 1475 1026
rect 1435 906 1475 909
rect 1437 900 1441 906
rect 1453 876 1457 880
rect 1423 872 1457 876
rect 1398 864 1402 872
rect 1445 864 1449 872
rect 1390 838 1394 844
rect 1406 838 1410 844
rect 1437 838 1441 844
rect 1453 838 1457 844
rect 1358 835 1413 838
rect 1358 742 1361 835
rect 1434 835 1463 838
rect 1394 787 1398 828
rect 1402 824 1445 828
rect 1412 803 1416 812
rect 1449 811 1453 828
rect 1442 807 1456 811
rect 1412 799 1422 803
rect 1472 803 1475 906
rect 1412 798 1416 799
rect 1449 787 1453 800
rect 1466 799 1475 803
rect 1394 783 1453 787
rect 1394 715 1398 783
rect 1407 773 1453 776
rect 1412 752 1416 762
rect 1449 760 1453 773
rect 1442 756 1456 760
rect 1412 748 1422 752
rect 1472 752 1475 799
rect 1412 742 1416 748
rect 1449 727 1453 749
rect 1466 748 1475 752
rect 771 631 783 635
rect 779 627 783 631
rect 683 624 726 627
rect 646 617 655 621
rect 544 605 639 609
rect 646 605 649 617
rect 683 613 687 624
rect 742 623 751 627
rect 779 623 787 627
rect 711 617 721 621
rect 675 609 687 613
rect 683 605 687 609
rect 646 601 655 605
rect 683 601 691 605
rect 717 598 721 617
rect 811 598 815 639
rect 532 594 815 598
rect 924 638 980 642
rect 988 709 1253 713
rect 1259 711 1398 715
rect 531 563 625 566
rect 531 531 535 545
rect 542 539 545 563
rect 621 560 625 563
rect 574 542 614 546
rect 574 539 578 542
rect 542 535 548 539
rect 574 535 581 539
rect 518 523 535 527
rect 542 523 545 535
rect 574 531 578 535
rect 610 531 614 542
rect 629 531 633 540
rect 568 527 578 531
rect 610 527 622 531
rect 629 527 670 531
rect 629 524 633 527
rect 471 518 496 521
rect 518 512 522 523
rect 542 519 548 523
rect 601 519 607 523
rect 351 508 522 512
rect 604 511 607 519
rect 621 511 625 514
rect 531 508 625 511
rect 351 504 355 508
rect 331 500 355 504
rect 331 484 335 500
rect 362 498 489 501
rect 531 499 648 502
rect 355 493 366 495
rect 355 491 362 493
rect 373 488 376 498
rect 471 495 475 498
rect 405 491 465 494
rect 405 488 408 491
rect 288 480 335 484
rect 346 481 358 485
rect 251 472 260 476
rect 231 468 244 472
rect 231 461 244 464
rect 192 460 244 461
rect 251 460 254 472
rect 288 468 292 480
rect 316 472 320 476
rect 280 464 292 468
rect 288 460 292 464
rect 192 457 235 460
rect 155 450 164 454
rect 53 438 148 442
rect 155 438 158 450
rect 192 446 196 457
rect 251 456 260 460
rect 288 456 296 460
rect 220 450 230 454
rect 184 442 196 446
rect 192 438 196 442
rect 155 434 164 438
rect 192 434 200 438
rect 226 431 230 450
rect 320 431 324 472
rect 331 460 335 480
rect 354 480 358 481
rect 362 480 366 488
rect 373 484 379 488
rect 404 484 411 488
rect 359 475 366 476
rect 354 472 366 475
rect 373 472 376 484
rect 404 480 408 484
rect 399 476 408 480
rect 373 468 379 472
rect 346 464 366 468
rect 331 456 366 460
rect 373 456 376 468
rect 404 464 408 476
rect 462 466 465 491
rect 527 487 535 491
rect 479 466 483 475
rect 399 460 408 464
rect 462 462 472 466
rect 479 462 498 466
rect 479 459 483 462
rect 331 436 335 456
rect 373 452 379 456
rect 451 452 457 456
rect 373 449 376 452
rect 454 446 457 452
rect 471 446 475 449
rect 494 447 498 462
rect 502 462 505 483
rect 531 478 535 487
rect 542 478 545 499
rect 630 496 634 499
rect 666 498 670 527
rect 678 511 836 514
rect 574 489 624 492
rect 574 486 577 489
rect 568 482 580 486
rect 542 474 548 478
rect 517 471 535 474
rect 512 470 535 471
rect 520 462 535 466
rect 542 462 545 474
rect 573 470 577 482
rect 568 466 577 470
rect 613 462 616 486
rect 621 467 624 489
rect 666 494 682 498
rect 661 486 682 490
rect 638 467 642 476
rect 651 478 682 482
rect 651 467 655 478
rect 621 463 631 467
rect 638 463 655 467
rect 663 470 682 474
rect 689 470 692 511
rect 780 505 812 508
rect 780 502 783 505
rect 775 498 783 502
rect 797 498 803 502
rect 779 494 783 498
rect 779 490 787 494
rect 779 478 783 490
rect 800 486 803 498
rect 797 482 803 486
rect 779 474 787 478
rect 800 470 803 482
rect 809 478 812 505
rect 818 507 822 511
rect 826 478 830 487
rect 809 474 819 478
rect 826 474 842 478
rect 826 471 830 474
rect 502 459 510 462
rect 507 451 510 459
rect 362 443 483 446
rect 520 435 524 462
rect 542 458 548 462
rect 610 458 616 462
rect 638 460 642 463
rect 613 447 616 458
rect 630 447 634 450
rect 531 444 642 447
rect 336 431 524 435
rect 663 437 667 470
rect 689 466 695 470
rect 797 466 803 470
rect 800 458 803 466
rect 818 458 822 461
rect 678 455 830 458
rect 708 442 802 445
rect 663 433 712 437
rect 663 431 667 433
rect 41 427 324 431
rect 536 427 667 431
rect 41 420 135 423
rect 52 396 55 420
rect 131 417 135 420
rect 536 419 540 427
rect 84 399 124 403
rect 84 396 88 399
rect 52 392 58 396
rect 84 392 91 396
rect 30 388 45 392
rect 22 380 45 384
rect 52 380 55 392
rect 84 388 88 392
rect 120 388 124 399
rect 139 388 143 397
rect 151 415 540 419
rect 151 388 155 415
rect 708 410 712 433
rect 719 418 722 442
rect 798 439 802 442
rect 751 421 795 425
rect 751 418 755 421
rect 719 414 725 418
rect 751 414 758 418
rect 511 407 686 410
rect 683 398 686 407
rect 700 403 712 406
rect 719 402 722 414
rect 751 410 755 414
rect 745 406 755 410
rect 791 410 795 421
rect 806 410 810 419
rect 838 418 842 474
rect 854 432 857 455
rect 791 406 799 410
rect 806 406 820 410
rect 806 403 810 406
rect 719 398 725 402
rect 778 398 784 402
rect 683 395 701 398
rect 78 384 88 388
rect 120 384 132 388
rect 139 384 155 388
rect 301 386 403 389
rect 426 387 553 390
rect 572 387 689 390
rect 139 381 143 384
rect 52 376 58 380
rect 111 376 117 380
rect 114 368 117 376
rect 131 368 135 371
rect 41 365 135 368
rect 278 363 282 369
rect 290 367 294 379
rect 301 367 304 386
rect 385 383 389 386
rect 333 378 379 381
rect 333 375 336 378
rect 327 371 339 375
rect 301 363 307 367
rect 278 359 294 363
rect 268 355 272 358
rect 268 351 294 355
rect 301 351 304 363
rect 332 359 336 371
rect 327 355 336 359
rect 301 347 307 351
rect 42 342 255 346
rect 259 343 294 347
rect 193 331 236 335
rect 156 324 165 328
rect 54 320 149 324
rect -703 308 11 312
rect -1186 299 -912 302
rect -1186 296 -1183 299
rect -916 296 -912 299
rect -1336 293 -1134 296
rect -1243 264 -1240 293
rect -1137 282 -1134 293
rect -916 293 -807 296
rect -1100 288 -964 292
rect -1137 278 -1128 282
rect -1206 274 -1144 278
rect -1243 260 -1234 264
rect -1351 256 -1250 260
rect -1336 238 -1316 242
rect -1330 232 -1326 238
rect -1322 205 -1318 212
rect -1305 205 -1302 247
rect -1351 201 -1329 205
rect -1322 201 -1302 205
rect -1295 205 -1291 256
rect -1280 238 -1266 242
rect -1279 232 -1275 238
rect -1271 205 -1267 212
rect -1254 209 -1250 252
rect -1243 248 -1240 260
rect -1206 256 -1202 274
rect -1172 264 -1169 270
rect -1178 260 -1169 264
rect -1214 252 -1202 256
rect -1206 248 -1202 252
rect -1243 244 -1234 248
rect -1206 244 -1198 248
rect -1243 241 -1240 244
rect -1172 242 -1169 260
rect -1137 266 -1134 278
rect -1100 274 -1096 288
rect -1072 278 -1070 282
rect -1108 270 -1096 274
rect -1100 266 -1096 270
rect -1144 259 -1141 266
rect -1137 262 -1128 266
rect -1100 262 -1092 266
rect -1137 256 -1134 262
rect -1062 251 -1058 288
rect -1144 247 -1058 251
rect -1206 227 -1160 231
rect -1243 217 -1240 220
rect -1243 213 -1234 217
rect -1295 201 -1278 205
rect -1271 201 -1250 205
rect -1243 201 -1240 213
rect -1206 209 -1202 227
rect -1172 217 -1169 219
rect -1178 213 -1169 217
rect -1214 205 -1202 209
rect -1206 201 -1202 205
rect -1322 198 -1318 201
rect -1271 198 -1267 201
rect -1243 197 -1234 201
rect -1206 197 -1198 201
rect -1243 191 -1240 197
rect -1330 182 -1326 188
rect -1279 182 -1275 188
rect -1172 182 -1169 213
rect -1164 205 -1160 227
rect -1144 213 -1140 247
rect -1137 217 -1134 223
rect -1137 213 -1128 217
rect -1164 201 -1144 205
rect -1137 201 -1134 213
rect -1100 209 -1096 239
rect -1052 217 -1049 278
rect -968 260 -964 288
rect -916 264 -913 293
rect -810 282 -807 293
rect -703 292 -699 308
rect -527 298 -253 301
rect -527 295 -524 298
rect -257 295 -253 298
rect -677 292 -475 295
rect -773 288 -699 292
rect -810 278 -801 282
rect -879 274 -817 278
rect -916 260 -907 264
rect -968 256 -923 260
rect -1008 238 -984 242
rect -1072 213 -1049 217
rect -1108 205 -1096 209
rect -1100 201 -1096 205
rect -1137 197 -1128 201
rect -1100 197 -1092 201
rect -1137 191 -1134 197
rect -1052 182 -1049 213
rect -1002 232 -998 238
rect -994 205 -990 212
rect -978 205 -973 247
rect -1013 201 -1001 205
rect -994 201 -973 205
rect -968 205 -964 256
rect -953 238 -939 242
rect -952 232 -948 238
rect -944 205 -940 212
rect -927 209 -923 252
rect -916 248 -913 260
rect -879 256 -875 274
rect -845 264 -842 270
rect -851 260 -842 264
rect -887 252 -875 256
rect -879 248 -875 252
rect -916 244 -907 248
rect -879 244 -871 248
rect -916 241 -913 244
rect -845 242 -842 260
rect -810 266 -807 278
rect -773 274 -769 288
rect -745 278 -743 282
rect -781 270 -769 274
rect -773 266 -769 270
rect -817 259 -814 266
rect -810 262 -801 266
rect -773 262 -765 266
rect -810 256 -807 262
rect -735 251 -731 288
rect -817 247 -731 251
rect -879 227 -833 231
rect -916 217 -913 220
rect -916 213 -907 217
rect -968 201 -951 205
rect -944 201 -923 205
rect -916 201 -913 213
rect -879 209 -875 227
rect -845 217 -842 219
rect -851 213 -842 217
rect -887 205 -875 209
rect -879 201 -875 205
rect -994 198 -990 201
rect -944 198 -940 201
rect -916 197 -907 201
rect -879 197 -871 201
rect -916 191 -913 197
rect -1002 182 -998 188
rect -952 182 -948 188
rect -845 182 -842 213
rect -837 205 -833 227
rect -817 213 -813 247
rect -810 217 -807 223
rect -810 213 -801 217
rect -837 201 -817 205
rect -810 201 -807 213
rect -773 209 -769 239
rect -725 217 -722 278
rect -584 263 -581 292
rect -478 281 -475 292
rect -257 292 -148 295
rect -441 287 -305 291
rect -478 277 -469 281
rect -547 273 -485 277
rect -584 259 -575 263
rect -692 255 -591 259
rect -677 237 -657 241
rect -745 213 -722 217
rect -781 205 -769 209
rect -773 201 -769 205
rect -810 197 -801 201
rect -773 197 -765 201
rect -810 191 -807 197
rect -725 182 -722 213
rect -671 231 -667 237
rect -663 204 -659 211
rect -646 204 -643 246
rect -692 200 -670 204
rect -663 200 -643 204
rect -636 204 -632 255
rect -621 237 -607 241
rect -620 231 -616 237
rect -612 204 -608 211
rect -595 208 -591 251
rect -584 247 -581 259
rect -547 255 -543 273
rect -513 263 -510 269
rect -519 259 -510 263
rect -555 251 -543 255
rect -547 247 -543 251
rect -584 243 -575 247
rect -547 243 -539 247
rect -584 240 -581 243
rect -513 241 -510 259
rect -478 265 -475 277
rect -441 273 -437 287
rect -413 277 -411 281
rect -449 269 -437 273
rect -441 265 -437 269
rect -485 258 -482 265
rect -478 261 -469 265
rect -441 261 -433 265
rect -478 255 -475 261
rect -403 250 -399 287
rect -485 246 -399 250
rect -547 226 -501 230
rect -584 216 -581 219
rect -584 212 -575 216
rect -636 200 -619 204
rect -612 200 -591 204
rect -584 200 -581 212
rect -547 208 -543 226
rect -513 216 -510 218
rect -519 212 -510 216
rect -555 204 -543 208
rect -547 200 -543 204
rect -663 197 -659 200
rect -612 197 -608 200
rect -1330 179 -722 182
rect -584 196 -575 200
rect -547 196 -539 200
rect -584 190 -581 196
rect -671 181 -667 187
rect -620 181 -616 187
rect -513 181 -510 212
rect -505 204 -501 226
rect -485 212 -481 246
rect -478 216 -475 222
rect -478 212 -469 216
rect -505 200 -485 204
rect -478 200 -475 212
rect -441 208 -437 238
rect -393 216 -390 277
rect -309 259 -305 287
rect -257 263 -254 292
rect -151 281 -148 292
rect -114 287 -40 291
rect -151 277 -142 281
rect -220 273 -158 277
rect -257 259 -248 263
rect -309 255 -264 259
rect -349 237 -325 241
rect -413 212 -390 216
rect -449 204 -437 208
rect -441 200 -437 204
rect -478 196 -469 200
rect -441 196 -433 200
rect -478 190 -475 196
rect -393 181 -390 212
rect -343 231 -339 237
rect -335 204 -331 211
rect -319 204 -314 246
rect -354 200 -342 204
rect -335 200 -314 204
rect -309 204 -305 255
rect -294 237 -280 241
rect -293 231 -289 237
rect -285 204 -281 211
rect -268 208 -264 251
rect -257 247 -254 259
rect -220 255 -216 273
rect -186 263 -183 269
rect -192 259 -183 263
rect -228 251 -216 255
rect -220 247 -216 251
rect -257 243 -248 247
rect -220 243 -212 247
rect -257 240 -254 243
rect -186 241 -183 259
rect -151 265 -148 277
rect -114 273 -110 287
rect -86 277 -84 281
rect -122 269 -110 273
rect -114 265 -110 269
rect -158 258 -155 265
rect -151 261 -142 265
rect -114 261 -106 265
rect -151 255 -148 261
rect -76 250 -72 287
rect -44 282 -40 287
rect 7 290 11 308
rect 54 290 58 320
rect 145 301 149 316
rect 156 312 159 324
rect 193 320 197 331
rect 221 324 224 328
rect 185 316 197 320
rect 193 312 197 316
rect 102 297 149 301
rect 65 290 74 294
rect 7 286 58 290
rect -44 278 14 282
rect -158 246 -72 250
rect -220 226 -174 230
rect -257 216 -254 219
rect -257 212 -248 216
rect -309 200 -292 204
rect -285 200 -264 204
rect -257 200 -254 212
rect -220 208 -216 226
rect -186 216 -183 218
rect -192 212 -183 216
rect -228 204 -216 208
rect -220 200 -216 204
rect -335 197 -331 200
rect -285 197 -281 200
rect -257 196 -248 200
rect -220 196 -212 200
rect -257 190 -254 196
rect -343 181 -339 187
rect -293 181 -289 187
rect -186 181 -183 212
rect -178 204 -174 226
rect -158 212 -154 246
rect -151 216 -148 222
rect -151 212 -142 216
rect -178 200 -158 204
rect -151 200 -148 212
rect -114 208 -110 238
rect -66 216 -63 277
rect -86 212 -63 216
rect -122 204 -110 208
rect -114 200 -110 204
rect -151 196 -142 200
rect -114 196 -106 200
rect -151 190 -148 196
rect -66 181 -63 212
rect 31 210 35 286
rect 47 278 58 282
rect 65 278 68 290
rect 102 286 106 297
rect 130 290 134 294
rect 94 282 106 286
rect 102 278 106 282
rect 54 260 58 278
rect 65 274 74 278
rect 102 274 110 278
rect 145 264 149 297
rect 156 308 165 312
rect 193 308 201 312
rect 156 299 160 308
rect 156 295 205 299
rect 156 272 160 295
rect 232 290 236 331
rect 251 299 255 342
rect 270 311 274 343
rect 282 335 294 339
rect 301 335 304 347
rect 332 343 336 355
rect 376 354 379 378
rect 427 377 430 382
rect 426 369 430 377
rect 437 377 440 387
rect 535 384 539 387
rect 469 380 529 383
rect 469 377 472 380
rect 437 373 443 377
rect 468 373 475 377
rect 393 354 397 363
rect 404 364 430 365
rect 409 361 430 364
rect 437 361 440 373
rect 468 369 472 373
rect 463 365 472 369
rect 437 357 443 361
rect 413 354 430 357
rect 376 350 386 354
rect 393 350 408 354
rect 393 347 397 350
rect 327 339 336 343
rect 282 308 286 335
rect 301 331 307 335
rect 364 334 367 335
rect 364 331 370 334
rect 367 325 370 331
rect 385 325 389 337
rect 290 322 389 325
rect 404 319 408 350
rect 418 353 430 354
rect 426 337 430 349
rect 437 345 440 357
rect 468 353 472 365
rect 526 355 529 380
rect 568 376 576 380
rect 572 366 576 376
rect 583 366 586 387
rect 671 384 675 387
rect 615 377 665 380
rect 615 374 618 377
rect 609 370 621 374
rect 543 355 547 364
rect 583 362 589 366
rect 559 358 576 362
rect 463 349 472 353
rect 526 351 536 355
rect 543 352 561 355
rect 543 351 548 352
rect 553 351 561 352
rect 543 348 547 351
rect 437 341 443 345
rect 515 344 518 345
rect 515 341 521 344
rect 437 338 440 341
rect 518 335 521 341
rect 535 335 539 338
rect 441 332 547 335
rect 557 321 561 351
rect 569 350 576 354
rect 583 350 586 362
rect 614 358 618 370
rect 609 354 618 358
rect 662 355 665 377
rect 698 379 701 395
rect 781 390 784 398
rect 798 390 802 393
rect 708 387 802 390
rect 816 384 820 406
rect 831 402 879 405
rect 876 390 879 402
rect 876 387 894 390
rect 711 380 820 384
rect 679 355 683 364
rect 711 357 715 380
rect 824 374 909 377
rect 718 366 894 369
rect 662 351 672 355
rect 679 351 688 355
rect 711 353 722 357
rect 569 341 573 350
rect 583 346 589 350
rect 620 346 621 350
rect 679 348 683 351
rect 620 335 623 346
rect 718 346 722 353
rect 711 338 722 342
rect 671 335 675 338
rect 599 332 683 335
rect 710 330 722 334
rect 582 323 681 327
rect 335 313 366 317
rect 404 315 461 319
rect 282 304 293 308
rect 289 302 293 304
rect 335 302 339 313
rect 582 309 586 323
rect 289 298 339 302
rect 347 305 586 309
rect 252 290 261 294
rect 232 286 245 290
rect 232 279 245 282
rect 193 278 245 279
rect 252 278 255 290
rect 289 286 293 298
rect 317 290 321 294
rect 347 294 351 305
rect 333 290 351 294
rect 281 282 293 286
rect 289 278 293 282
rect 193 275 236 278
rect 156 268 165 272
rect 54 256 149 260
rect 156 256 159 268
rect 193 264 197 275
rect 252 274 261 278
rect 289 274 297 278
rect 221 268 231 272
rect 185 260 197 264
rect 193 256 197 260
rect 156 252 165 256
rect 193 252 201 256
rect 227 249 231 268
rect 289 264 293 274
rect 262 258 288 262
rect 321 249 325 290
rect 42 245 325 249
rect 333 241 337 290
rect 365 273 578 277
rect 516 262 559 266
rect 479 255 488 259
rect 42 238 136 241
rect 53 214 56 238
rect 132 235 136 238
rect 153 237 337 241
rect 377 251 472 255
rect 85 217 125 221
rect 85 214 89 217
rect 53 210 59 214
rect 85 210 92 214
rect 31 206 46 210
rect 23 198 46 202
rect 53 198 56 210
rect 85 206 89 210
rect 121 206 125 217
rect 140 206 144 215
rect 153 206 157 237
rect 79 202 89 206
rect 121 202 133 206
rect 140 202 157 206
rect 140 199 144 202
rect 53 194 59 198
rect 112 194 118 198
rect 115 186 118 194
rect 132 186 136 189
rect 42 183 136 186
rect -671 178 -63 181
rect 258 174 261 229
rect 270 190 274 227
rect 317 225 369 229
rect 365 221 369 225
rect 377 221 381 251
rect 468 232 472 247
rect 479 243 482 255
rect 516 251 520 262
rect 544 255 547 259
rect 508 247 520 251
rect 516 243 520 247
rect 425 228 472 232
rect 388 221 397 225
rect 365 217 381 221
rect 336 213 341 214
rect 336 209 381 213
rect 388 209 391 221
rect 425 217 429 228
rect 453 221 457 225
rect 417 213 429 217
rect 425 209 429 213
rect 285 201 348 204
rect 270 187 339 190
rect 270 186 274 187
rect 258 171 327 174
rect 43 159 256 163
rect 194 148 237 152
rect 157 141 166 145
rect 55 137 150 141
rect -703 120 11 124
rect -1186 112 -912 115
rect -1186 109 -1183 112
rect -916 109 -912 112
rect -1336 106 -1134 109
rect -1243 77 -1240 106
rect -1137 95 -1134 106
rect -916 106 -807 109
rect -1100 101 -964 105
rect -1137 91 -1128 95
rect -1206 87 -1144 91
rect -1243 73 -1234 77
rect -1351 69 -1250 73
rect -1336 51 -1316 55
rect -1330 45 -1326 51
rect -1322 18 -1318 25
rect -1305 18 -1302 60
rect -1351 14 -1329 18
rect -1322 14 -1302 18
rect -1295 18 -1291 69
rect -1280 51 -1266 55
rect -1279 45 -1275 51
rect -1271 18 -1267 25
rect -1254 22 -1250 65
rect -1243 61 -1240 73
rect -1206 69 -1202 87
rect -1172 77 -1169 83
rect -1178 73 -1169 77
rect -1214 65 -1202 69
rect -1206 61 -1202 65
rect -1243 57 -1234 61
rect -1206 57 -1198 61
rect -1243 54 -1240 57
rect -1172 55 -1169 73
rect -1137 79 -1134 91
rect -1100 87 -1096 101
rect -1072 91 -1070 95
rect -1108 83 -1096 87
rect -1100 79 -1096 83
rect -1144 72 -1141 79
rect -1137 75 -1128 79
rect -1100 75 -1092 79
rect -1137 69 -1134 75
rect -1062 64 -1058 101
rect -1144 60 -1058 64
rect -1206 40 -1160 44
rect -1243 30 -1240 33
rect -1243 26 -1234 30
rect -1295 14 -1278 18
rect -1271 14 -1250 18
rect -1243 14 -1240 26
rect -1206 22 -1202 40
rect -1172 30 -1169 32
rect -1178 26 -1169 30
rect -1214 18 -1202 22
rect -1206 14 -1202 18
rect -1322 11 -1318 14
rect -1271 11 -1267 14
rect -1243 10 -1234 14
rect -1206 10 -1198 14
rect -1243 4 -1240 10
rect -1330 -5 -1326 1
rect -1279 -5 -1275 1
rect -1172 -5 -1169 26
rect -1164 18 -1160 40
rect -1144 26 -1140 60
rect -1137 30 -1134 36
rect -1137 26 -1128 30
rect -1164 14 -1144 18
rect -1137 14 -1134 26
rect -1100 22 -1096 52
rect -1052 30 -1049 91
rect -968 73 -964 101
rect -916 77 -913 106
rect -810 95 -807 106
rect -703 105 -699 120
rect -527 111 -253 114
rect -527 108 -524 111
rect -257 108 -253 111
rect -677 105 -475 108
rect -773 101 -699 105
rect -810 91 -801 95
rect -879 87 -817 91
rect -916 73 -907 77
rect -968 69 -923 73
rect -1008 51 -984 55
rect -1072 26 -1049 30
rect -1108 18 -1096 22
rect -1100 14 -1096 18
rect -1137 10 -1128 14
rect -1100 10 -1092 14
rect -1137 4 -1134 10
rect -1052 -5 -1049 26
rect -1002 45 -998 51
rect -994 18 -990 25
rect -978 18 -973 60
rect -1013 14 -1001 18
rect -994 14 -973 18
rect -968 18 -964 69
rect -953 51 -939 55
rect -952 45 -948 51
rect -944 18 -940 25
rect -927 22 -923 65
rect -916 61 -913 73
rect -879 69 -875 87
rect -845 77 -842 83
rect -851 73 -842 77
rect -887 65 -875 69
rect -879 61 -875 65
rect -916 57 -907 61
rect -879 57 -871 61
rect -916 54 -913 57
rect -845 55 -842 73
rect -810 79 -807 91
rect -773 87 -769 101
rect -745 91 -743 95
rect -781 83 -769 87
rect -773 79 -769 83
rect -817 72 -814 79
rect -810 75 -801 79
rect -773 75 -765 79
rect -810 69 -807 75
rect -735 64 -731 101
rect -817 60 -731 64
rect -879 40 -833 44
rect -916 30 -913 33
rect -916 26 -907 30
rect -968 14 -951 18
rect -944 14 -923 18
rect -916 14 -913 26
rect -879 22 -875 40
rect -845 30 -842 32
rect -851 26 -842 30
rect -887 18 -875 22
rect -879 14 -875 18
rect -994 11 -990 14
rect -944 11 -940 14
rect -916 10 -907 14
rect -879 10 -871 14
rect -916 4 -913 10
rect -1002 -5 -998 1
rect -952 -5 -948 1
rect -845 -5 -842 26
rect -837 18 -833 40
rect -817 26 -813 60
rect -810 30 -807 36
rect -810 26 -801 30
rect -837 14 -817 18
rect -810 14 -807 26
rect -773 22 -769 52
rect -725 30 -722 91
rect -584 76 -581 105
rect -478 94 -475 105
rect -257 105 -148 108
rect -441 100 -305 104
rect -478 90 -469 94
rect -547 86 -485 90
rect -584 72 -575 76
rect -692 68 -591 72
rect -677 50 -657 54
rect -745 26 -722 30
rect -781 18 -769 22
rect -773 14 -769 18
rect -810 10 -801 14
rect -773 10 -765 14
rect -810 4 -807 10
rect -725 -5 -722 26
rect -671 44 -667 50
rect -663 17 -659 24
rect -646 17 -643 59
rect -692 13 -670 17
rect -663 13 -643 17
rect -636 17 -632 68
rect -621 50 -607 54
rect -620 44 -616 50
rect -612 17 -608 24
rect -595 21 -591 64
rect -584 60 -581 72
rect -547 68 -543 86
rect -513 76 -510 82
rect -519 72 -510 76
rect -555 64 -543 68
rect -547 60 -543 64
rect -584 56 -575 60
rect -547 56 -539 60
rect -584 53 -581 56
rect -513 54 -510 72
rect -478 78 -475 90
rect -441 86 -437 100
rect -413 90 -411 94
rect -449 82 -437 86
rect -441 78 -437 82
rect -485 71 -482 78
rect -478 74 -469 78
rect -441 74 -433 78
rect -478 68 -475 74
rect -403 63 -399 100
rect -485 59 -399 63
rect -547 39 -501 43
rect -584 29 -581 32
rect -584 25 -575 29
rect -636 13 -619 17
rect -612 13 -591 17
rect -584 13 -581 25
rect -547 21 -543 39
rect -513 29 -510 31
rect -519 25 -510 29
rect -555 17 -543 21
rect -547 13 -543 17
rect -663 10 -659 13
rect -612 10 -608 13
rect -1330 -8 -722 -5
rect -584 9 -575 13
rect -547 9 -539 13
rect -584 3 -581 9
rect -671 -6 -667 0
rect -620 -6 -616 0
rect -513 -6 -510 25
rect -505 17 -501 39
rect -485 25 -481 59
rect -478 29 -475 35
rect -478 25 -469 29
rect -505 13 -485 17
rect -478 13 -475 25
rect -441 21 -437 51
rect -393 29 -390 90
rect -309 72 -305 100
rect -257 76 -254 105
rect -151 94 -148 105
rect 7 107 11 120
rect 55 107 59 137
rect 146 118 150 133
rect 157 129 160 141
rect 194 137 198 148
rect 222 141 225 145
rect 186 133 198 137
rect 194 129 198 133
rect 103 114 150 118
rect 66 107 75 111
rect -114 100 -40 104
rect 7 103 59 107
rect -151 90 -142 94
rect -220 86 -158 90
rect -257 72 -248 76
rect -309 68 -264 72
rect -349 50 -325 54
rect -413 25 -390 29
rect -449 17 -437 21
rect -441 13 -437 17
rect -478 9 -469 13
rect -441 9 -433 13
rect -478 3 -475 9
rect -393 -6 -390 25
rect -343 44 -339 50
rect -335 17 -331 24
rect -319 17 -314 59
rect -354 13 -342 17
rect -335 13 -314 17
rect -309 17 -305 68
rect -294 50 -280 54
rect -293 44 -289 50
rect -285 17 -281 24
rect -268 21 -264 64
rect -257 60 -254 72
rect -220 68 -216 86
rect -186 76 -183 82
rect -192 72 -183 76
rect -228 64 -216 68
rect -220 60 -216 64
rect -257 56 -248 60
rect -220 56 -212 60
rect -257 53 -254 56
rect -186 54 -183 72
rect -151 78 -148 90
rect -114 86 -110 100
rect -86 90 -84 94
rect -122 82 -110 86
rect -114 78 -110 82
rect -158 71 -155 78
rect -151 74 -142 78
rect -114 74 -106 78
rect -151 68 -148 74
rect -76 63 -72 100
rect -44 99 -40 100
rect -44 95 15 99
rect -158 59 -72 63
rect -220 39 -174 43
rect -257 29 -254 32
rect -257 25 -248 29
rect -309 13 -292 17
rect -285 13 -264 17
rect -257 13 -254 25
rect -220 21 -216 39
rect -186 29 -183 31
rect -192 25 -183 29
rect -228 17 -216 21
rect -220 13 -216 17
rect -335 10 -331 13
rect -285 10 -281 13
rect -257 9 -248 13
rect -220 9 -212 13
rect -257 3 -254 9
rect -343 -6 -339 0
rect -293 -6 -289 0
rect -186 -6 -183 25
rect -178 17 -174 39
rect -158 25 -154 59
rect -151 29 -148 35
rect -151 25 -142 29
rect -178 13 -158 17
rect -151 13 -148 25
rect -114 21 -110 51
rect -66 29 -63 90
rect -86 25 -63 29
rect -122 17 -110 21
rect -114 13 -110 17
rect -151 9 -142 13
rect -114 9 -106 13
rect -151 3 -148 9
rect -66 -6 -63 25
rect 32 27 36 103
rect 48 95 59 99
rect 66 95 69 107
rect 103 103 107 114
rect 131 107 135 111
rect 95 99 107 103
rect 103 95 107 99
rect 55 77 59 95
rect 66 91 75 95
rect 103 91 111 95
rect 146 81 150 114
rect 157 125 166 129
rect 194 125 202 129
rect 157 116 161 125
rect 157 112 206 116
rect 157 89 161 112
rect 233 107 237 148
rect 252 116 256 159
rect 324 120 327 171
rect 336 136 339 187
rect 324 117 333 120
rect 253 107 262 111
rect 233 103 246 107
rect 233 96 246 99
rect 194 95 246 96
rect 253 95 256 107
rect 290 103 294 115
rect 318 107 322 111
rect 282 99 294 103
rect 290 95 294 99
rect 194 92 237 95
rect 157 85 166 89
rect 55 73 150 77
rect 157 73 160 85
rect 194 81 198 92
rect 253 91 262 95
rect 290 91 298 95
rect 222 85 232 89
rect 186 77 198 81
rect 194 73 198 77
rect 157 69 166 73
rect 194 69 202 73
rect 228 66 232 85
rect 290 81 294 91
rect 290 77 304 81
rect 322 66 326 107
rect 330 99 333 117
rect 345 115 348 201
rect 377 191 381 209
rect 388 205 397 209
rect 425 205 433 209
rect 468 195 472 228
rect 479 239 488 243
rect 516 239 524 243
rect 479 230 483 239
rect 479 226 528 230
rect 479 203 483 226
rect 555 221 559 262
rect 574 230 578 273
rect 657 247 661 323
rect 677 303 681 323
rect 709 322 722 326
rect 709 313 713 322
rect 702 309 713 313
rect 718 303 722 318
rect 729 314 732 366
rect 876 363 880 366
rect 841 357 870 360
rect 841 354 844 357
rect 835 350 847 354
rect 840 338 844 350
rect 860 346 863 354
rect 857 342 863 346
rect 840 334 847 338
rect 840 322 844 334
rect 860 330 863 342
rect 867 334 870 357
rect 884 334 888 343
rect 867 330 877 334
rect 884 330 895 334
rect 857 326 863 330
rect 884 327 888 330
rect 840 318 847 322
rect 860 314 863 326
rect 729 310 735 314
rect 857 313 863 314
rect 876 313 880 317
rect 857 310 880 313
rect 729 304 732 310
rect 677 299 722 303
rect 860 300 863 310
rect 741 297 863 300
rect 906 293 909 374
rect 681 290 909 293
rect 657 243 667 247
rect 612 229 670 233
rect 575 221 584 225
rect 555 217 568 221
rect 555 210 568 213
rect 516 209 568 210
rect 575 209 578 221
rect 612 217 616 229
rect 640 221 644 225
rect 604 213 616 217
rect 612 209 616 213
rect 516 206 559 209
rect 479 199 488 203
rect 377 187 472 191
rect 479 187 482 199
rect 516 195 520 206
rect 575 205 584 209
rect 612 205 620 209
rect 544 199 554 203
rect 508 191 520 195
rect 516 187 520 191
rect 479 183 488 187
rect 516 183 524 187
rect 550 180 554 199
rect 644 180 648 221
rect 681 202 684 290
rect 924 278 928 638
rect 988 629 992 709
rect 1259 703 1263 711
rect 937 625 992 629
rect 999 699 1263 703
rect 937 290 941 625
rect 999 616 1003 699
rect 951 612 1003 616
rect 951 301 955 612
rect 951 297 1251 301
rect 937 286 1241 290
rect 787 274 928 278
rect 787 233 791 274
rect 990 270 1203 274
rect 1141 259 1184 263
rect 835 242 929 245
rect 697 230 791 233
rect 696 229 791 230
rect 689 219 806 222
rect 681 198 693 202
rect 700 198 703 219
rect 788 216 792 219
rect 732 209 782 212
rect 732 206 735 209
rect 726 202 738 206
rect 700 194 706 198
rect 678 190 693 194
rect 365 176 648 180
rect 689 179 693 186
rect 700 182 703 194
rect 731 190 735 202
rect 726 186 735 190
rect 771 182 774 206
rect 779 187 782 209
rect 813 214 817 242
rect 846 218 849 242
rect 925 239 929 242
rect 878 221 918 225
rect 878 218 882 221
rect 846 214 852 218
rect 878 214 885 218
rect 813 210 839 214
rect 816 205 839 206
rect 821 202 839 205
rect 846 202 849 214
rect 878 210 882 214
rect 914 210 918 221
rect 933 210 937 219
rect 990 218 994 254
rect 1104 252 1113 256
rect 1002 248 1097 252
rect 1002 218 1006 248
rect 1093 229 1097 244
rect 1104 240 1107 252
rect 1141 248 1145 259
rect 1169 252 1172 256
rect 1133 244 1145 248
rect 1141 240 1145 244
rect 1050 225 1097 229
rect 1013 218 1022 222
rect 990 214 1006 218
rect 872 206 882 210
rect 914 206 926 210
rect 933 206 954 210
rect 933 203 937 206
rect 846 198 852 202
rect 905 198 911 202
rect 796 187 800 196
rect 908 190 911 198
rect 925 190 929 193
rect 835 187 929 190
rect 779 183 789 187
rect 796 183 828 187
rect 669 176 693 179
rect 700 178 706 182
rect 768 178 774 182
rect 796 180 800 183
rect 771 167 774 178
rect 788 167 792 170
rect 712 164 800 167
rect 382 150 474 154
rect 364 135 375 139
rect 371 127 375 135
rect 382 135 386 150
rect 405 138 467 142
rect 405 135 409 138
rect 382 131 389 135
rect 405 131 413 135
rect 361 123 365 127
rect 361 119 375 123
rect 382 119 386 131
rect 405 127 409 131
rect 399 123 409 127
rect 382 115 389 119
rect 345 111 375 115
rect 341 105 375 107
rect 336 103 375 105
rect 382 103 386 115
rect 405 111 409 123
rect 399 107 409 111
rect 463 107 467 138
rect 470 136 474 150
rect 508 148 606 151
rect 509 138 512 143
rect 508 129 512 138
rect 519 129 522 148
rect 603 145 607 148
rect 551 140 600 143
rect 551 137 554 140
rect 545 133 557 137
rect 519 125 525 129
rect 499 121 512 125
rect 382 99 389 103
rect 330 95 375 99
rect 337 89 375 91
rect 342 87 375 89
rect 382 87 386 99
rect 405 95 409 107
rect 463 103 471 107
rect 478 100 482 116
rect 494 113 512 117
rect 519 113 522 125
rect 550 121 554 133
rect 545 117 554 121
rect 494 112 499 113
rect 399 91 409 95
rect 470 87 474 90
rect 382 83 389 87
rect 443 84 474 87
rect 504 98 507 108
rect 519 109 525 113
rect 443 83 446 84
rect 382 77 386 83
rect 43 62 326 66
rect 43 55 137 58
rect 478 56 482 90
rect 513 89 516 97
rect 519 97 522 109
rect 550 105 554 117
rect 597 116 600 140
rect 636 139 763 142
rect 824 139 828 183
rect 950 181 954 206
rect 980 206 1006 210
rect 1013 206 1016 218
rect 1050 214 1054 225
rect 1078 218 1082 222
rect 1042 210 1054 214
rect 1050 206 1054 210
rect 1002 188 1006 206
rect 1013 202 1022 206
rect 1050 202 1058 206
rect 1093 192 1097 225
rect 1104 236 1113 240
rect 1141 236 1149 240
rect 1104 227 1108 236
rect 1104 223 1153 227
rect 1104 200 1108 223
rect 1180 218 1184 259
rect 1199 227 1203 270
rect 1200 218 1209 222
rect 1180 214 1193 218
rect 1180 207 1193 210
rect 1141 206 1193 207
rect 1200 206 1203 218
rect 1237 214 1241 286
rect 1247 236 1251 297
rect 1247 232 1283 236
rect 1265 218 1269 222
rect 1229 210 1241 214
rect 1237 206 1241 210
rect 1141 203 1184 206
rect 1104 196 1113 200
rect 1002 184 1097 188
rect 1104 184 1107 196
rect 1141 192 1145 203
rect 1200 202 1209 206
rect 1237 202 1245 206
rect 1169 196 1179 200
rect 1133 188 1145 192
rect 1141 184 1145 188
rect 844 177 954 181
rect 1104 180 1113 184
rect 1141 180 1149 184
rect 1175 177 1179 196
rect 1269 177 1273 218
rect 647 129 650 139
rect 745 136 749 139
rect 824 136 835 139
rect 679 132 739 135
rect 679 129 682 132
rect 597 112 604 116
rect 611 109 615 125
rect 637 124 640 129
rect 647 125 653 129
rect 678 125 685 129
rect 636 121 640 124
rect 625 115 640 117
rect 630 113 640 115
rect 647 113 650 125
rect 678 121 682 125
rect 673 117 682 121
rect 647 109 653 113
rect 545 101 554 105
rect 519 93 525 97
rect 582 93 588 97
rect 585 87 588 93
rect 603 87 607 99
rect 534 84 607 87
rect 636 107 640 109
rect 611 75 615 99
rect 624 104 640 107
rect 624 103 629 104
rect 647 97 650 109
rect 678 105 682 117
rect 736 107 739 132
rect 831 133 835 136
rect 844 129 848 177
rect 990 173 1273 177
rect 1279 167 1283 232
rect 1059 163 1283 167
rect 856 145 1031 149
rect 844 125 849 129
rect 753 107 757 116
rect 770 117 849 121
rect 770 107 774 117
rect 673 101 682 105
rect 736 103 746 107
rect 753 103 774 107
rect 787 109 849 113
rect 753 100 757 103
rect 647 93 653 97
rect 725 93 731 97
rect 647 90 650 93
rect 728 87 731 93
rect 745 87 749 90
rect 636 84 757 87
rect 787 75 791 109
rect 611 71 791 75
rect 799 101 849 105
rect 799 56 803 101
rect 837 93 849 97
rect 845 83 849 89
rect 856 85 860 145
rect 987 137 1024 141
rect 1028 140 1031 145
rect 1028 137 1038 140
rect 987 133 991 137
rect 984 129 991 133
rect 1006 129 1013 133
rect 987 125 991 129
rect 987 121 996 125
rect 987 109 991 121
rect 1009 117 1013 129
rect 1006 113 1013 117
rect 987 105 996 109
rect 987 93 991 105
rect 1009 101 1013 113
rect 1020 105 1024 137
rect 1034 134 1038 137
rect 1042 105 1046 114
rect 1059 105 1063 163
rect 1020 101 1035 105
rect 1042 101 1063 105
rect 1006 97 1013 101
rect 1042 98 1046 101
rect 987 89 996 93
rect 1009 86 1013 97
rect 1034 86 1038 88
rect 1009 85 1038 86
rect 54 31 57 55
rect 133 52 137 55
rect 156 52 440 56
rect 478 52 803 56
rect 813 79 849 83
rect 856 81 864 85
rect 1006 82 1038 85
rect 1006 81 1013 82
rect 86 34 126 38
rect 86 31 90 34
rect 54 27 60 31
rect 86 27 93 31
rect 32 23 47 27
rect 24 15 47 19
rect 54 15 57 27
rect 86 23 90 27
rect 122 23 126 34
rect 141 23 145 32
rect 156 23 160 52
rect 436 47 440 52
rect 813 47 817 79
rect 436 43 817 47
rect 80 19 90 23
rect 122 19 134 23
rect 141 19 160 23
rect 141 16 145 19
rect 54 11 60 15
rect 113 11 119 15
rect 116 3 119 11
rect 133 3 137 6
rect 43 0 137 3
rect -671 -9 -63 -6
<< metal2 >>
rect 655 1340 658 1352
rect 797 1340 800 1352
rect 937 1340 940 1352
rect 1082 1340 1085 1352
rect 1227 1340 1230 1352
rect 1372 1340 1375 1352
rect 683 1305 693 1309
rect 825 1305 835 1309
rect 965 1305 975 1309
rect 1110 1305 1120 1309
rect 1255 1305 1265 1309
rect 1400 1305 1410 1309
rect 680 1264 683 1304
rect 710 1255 713 1268
rect 822 1264 825 1304
rect 649 1252 713 1255
rect 852 1255 855 1268
rect 962 1264 965 1304
rect 791 1252 855 1255
rect 992 1255 995 1268
rect 1107 1264 1110 1304
rect 931 1252 995 1255
rect 1137 1255 1140 1268
rect 1252 1264 1255 1304
rect 1076 1252 1140 1255
rect 1282 1255 1285 1268
rect 1397 1264 1400 1304
rect 1221 1252 1285 1255
rect 1427 1255 1430 1268
rect 1366 1252 1430 1255
rect 700 1233 713 1236
rect 842 1233 855 1236
rect 982 1233 995 1236
rect 1127 1233 1140 1236
rect 1272 1233 1285 1236
rect 1417 1233 1430 1236
rect -611 1155 -354 1158
rect 701 1161 712 1164
rect -611 1103 -608 1155
rect -641 1100 -599 1103
rect -651 1091 -625 1094
rect -601 1090 -585 1093
rect -585 1077 -580 1088
rect -512 1076 -509 1089
rect -493 1079 -490 1140
rect -405 1131 -393 1134
rect -481 1106 -441 1109
rect -440 1096 -436 1106
rect -493 1076 -477 1079
rect -357 1057 -354 1155
rect -335 1123 -261 1126
rect -335 1099 -332 1123
rect -313 1100 -272 1103
rect -274 1090 -258 1093
rect -257 1077 -254 1088
rect -185 1076 -182 1089
rect -166 1079 -163 1140
rect -78 1131 -66 1134
rect -154 1106 -114 1109
rect -113 1096 -109 1106
rect 663 1086 666 1157
rect 686 1105 689 1146
rect 696 1144 699 1160
rect 843 1161 854 1164
rect 663 1083 690 1086
rect 805 1086 808 1157
rect 828 1105 831 1146
rect 838 1144 841 1160
rect 983 1161 994 1164
rect 805 1083 832 1086
rect 945 1086 948 1157
rect 968 1105 971 1146
rect 978 1144 981 1160
rect 1128 1161 1139 1164
rect 945 1083 972 1086
rect 1090 1086 1093 1157
rect 1113 1105 1116 1146
rect 1123 1144 1126 1160
rect 1273 1161 1284 1164
rect 1090 1083 1117 1086
rect 1235 1086 1238 1157
rect 1258 1105 1261 1146
rect 1268 1144 1271 1160
rect 1418 1161 1429 1164
rect 1235 1083 1262 1086
rect 1380 1086 1383 1157
rect 1403 1105 1406 1146
rect 1413 1144 1416 1160
rect 1380 1083 1407 1086
rect -166 1076 -150 1079
rect 631 1061 732 1064
rect 316 1003 319 1041
rect 477 1020 480 1027
rect 477 1017 576 1020
rect 477 1011 480 1017
rect 449 1008 480 1011
rect -1271 995 -1014 998
rect -1271 943 -1268 995
rect -1301 940 -1259 943
rect -1311 931 -1285 934
rect -1261 930 -1245 933
rect -1245 917 -1240 928
rect -1172 916 -1169 929
rect -1153 919 -1150 980
rect -1065 971 -1053 974
rect -1141 946 -1101 949
rect -1100 936 -1096 946
rect -1153 916 -1137 919
rect -1017 897 -1014 995
rect -612 991 -355 994
rect 449 997 452 1008
rect 461 1000 501 1003
rect 573 999 576 1017
rect 390 994 452 997
rect -995 963 -921 966
rect -995 939 -992 963
rect -973 940 -932 943
rect -934 930 -918 933
rect -917 917 -914 928
rect -845 916 -842 929
rect -826 919 -823 980
rect -738 971 -726 974
rect -814 946 -774 949
rect -773 936 -769 946
rect -612 939 -609 991
rect -642 936 -600 939
rect -652 927 -626 930
rect -602 926 -586 929
rect -826 916 -810 919
rect -586 913 -581 924
rect -513 912 -510 925
rect -494 915 -491 976
rect -406 967 -394 970
rect -482 942 -442 945
rect -441 932 -437 942
rect -494 912 -478 915
rect -358 893 -355 991
rect -336 959 -262 962
rect -336 935 -333 959
rect -314 936 -273 939
rect -275 926 -259 929
rect -258 913 -255 924
rect -186 912 -183 925
rect -167 915 -164 976
rect -79 967 -67 970
rect -155 942 -115 945
rect -114 932 -110 942
rect -167 912 -151 915
rect 65 915 68 953
rect 285 947 289 968
rect 285 943 339 947
rect 226 932 229 939
rect 241 932 325 935
rect 226 929 244 932
rect 226 923 229 929
rect 198 920 229 923
rect 198 909 201 920
rect 210 912 250 915
rect 322 911 325 932
rect 335 925 339 943
rect 139 906 201 909
rect 19 894 42 898
rect 23 823 27 894
rect -1271 756 -1014 759
rect -1271 704 -1268 756
rect -1301 701 -1259 704
rect -1311 692 -1285 695
rect -1261 691 -1245 694
rect -1245 678 -1240 689
rect -1172 677 -1169 690
rect -1153 680 -1150 741
rect -1065 732 -1053 735
rect -1141 707 -1101 710
rect -1100 697 -1096 707
rect -1153 677 -1137 680
rect -1017 658 -1014 756
rect -612 755 -355 758
rect -995 724 -921 727
rect -995 700 -992 724
rect -973 701 -932 704
rect -934 691 -918 694
rect -917 678 -914 689
rect -845 677 -842 690
rect -826 680 -823 741
rect -738 732 -726 735
rect -814 707 -774 710
rect -773 697 -769 707
rect -612 703 -609 755
rect -642 700 -600 703
rect -652 691 -626 694
rect -602 690 -586 693
rect -826 677 -810 680
rect -586 677 -581 688
rect -513 676 -510 689
rect -494 679 -491 740
rect -406 731 -394 734
rect -482 706 -442 709
rect -441 696 -437 706
rect -494 676 -478 679
rect -358 657 -355 755
rect -336 723 -262 726
rect -336 699 -333 723
rect -314 700 -273 703
rect -275 690 -259 693
rect -258 677 -255 688
rect -186 676 -183 689
rect -167 679 -164 740
rect 64 735 67 773
rect 225 752 228 759
rect 225 749 324 752
rect 225 743 228 749
rect 197 740 228 743
rect -79 731 -67 734
rect 197 729 200 740
rect 209 732 249 735
rect 321 731 324 749
rect 335 748 339 865
rect 330 744 339 748
rect 138 726 200 729
rect 18 714 41 718
rect 330 717 334 744
rect -155 706 -115 709
rect -114 696 -110 706
rect -167 676 -151 679
rect 22 643 26 714
rect 345 703 348 892
rect 447 761 450 846
rect 631 810 634 1061
rect 773 1061 874 1064
rect 655 1013 658 1025
rect 683 978 693 982
rect 680 937 683 977
rect 710 928 713 941
rect 649 925 713 928
rect 700 906 713 909
rect 701 833 712 838
rect 686 810 689 819
rect 696 817 699 833
rect 631 807 689 810
rect 773 810 776 1061
rect 913 1061 1014 1064
rect 797 1013 800 1025
rect 825 978 835 982
rect 822 937 825 977
rect 852 928 855 941
rect 791 925 855 928
rect 842 906 855 909
rect 843 833 854 838
rect 828 810 831 819
rect 838 817 841 833
rect 773 807 831 810
rect 913 810 916 1061
rect 1058 1061 1159 1064
rect 937 1013 940 1025
rect 965 978 975 982
rect 962 937 965 977
rect 992 928 995 941
rect 931 925 995 928
rect 982 906 995 909
rect 983 833 994 838
rect 968 810 971 819
rect 978 817 981 833
rect 913 807 971 810
rect 1058 810 1061 1061
rect 1203 1061 1304 1064
rect 1082 1013 1085 1025
rect 1110 978 1120 982
rect 1107 937 1110 977
rect 1137 928 1140 941
rect 1076 925 1140 928
rect 1127 906 1140 909
rect 1128 833 1139 838
rect 1113 810 1116 819
rect 1123 817 1126 833
rect 1058 807 1116 810
rect 1203 810 1206 1061
rect 1348 1061 1449 1064
rect 1227 1013 1230 1025
rect 1255 978 1265 982
rect 1252 937 1255 977
rect 1282 928 1285 941
rect 1221 925 1285 928
rect 1272 906 1285 909
rect 1273 833 1284 838
rect 1258 810 1261 819
rect 1268 817 1271 833
rect 1203 807 1261 810
rect 1348 810 1351 1061
rect 1372 1013 1375 1025
rect 1400 978 1410 982
rect 1397 937 1400 977
rect 1427 928 1430 941
rect 1366 925 1430 928
rect 1417 906 1430 909
rect 1418 833 1429 838
rect 1403 810 1406 819
rect 1413 817 1416 833
rect 1348 807 1406 810
rect 538 788 556 791
rect 380 758 450 761
rect 380 724 383 758
rect 553 742 556 788
rect 686 777 689 807
rect 695 767 698 793
rect 828 777 831 807
rect 837 767 840 793
rect 968 777 971 807
rect 977 767 980 793
rect 1113 777 1116 807
rect 1122 767 1125 793
rect 1258 777 1261 807
rect 1267 767 1270 793
rect 1403 777 1406 807
rect 1412 767 1415 793
rect 513 739 556 742
rect 380 721 483 724
rect 444 702 446 707
rect 289 666 292 692
rect 168 663 292 666
rect 168 615 171 663
rect 345 656 348 698
rect 253 653 348 656
rect 157 612 171 615
rect -1271 542 -1014 545
rect -1271 490 -1268 542
rect -1301 487 -1259 490
rect -1311 478 -1285 481
rect -1261 477 -1245 480
rect -1245 464 -1240 475
rect -1172 463 -1169 476
rect -1153 466 -1150 527
rect -1065 518 -1053 521
rect -1141 493 -1101 496
rect -1100 483 -1096 493
rect -1153 463 -1137 466
rect -1017 444 -1014 542
rect -612 541 -355 544
rect -995 510 -921 513
rect -995 486 -992 510
rect -973 487 -932 490
rect -934 477 -918 480
rect -917 464 -914 475
rect -845 463 -842 476
rect -826 466 -823 527
rect -738 518 -726 521
rect -814 493 -774 496
rect -773 483 -769 493
rect -612 489 -609 541
rect -642 486 -600 489
rect -652 477 -626 480
rect -602 476 -586 479
rect -826 463 -810 466
rect -586 463 -581 474
rect -513 462 -510 475
rect -494 465 -491 526
rect -406 517 -394 520
rect -482 492 -442 495
rect -441 482 -437 492
rect -494 462 -478 465
rect -358 443 -355 541
rect 157 530 160 612
rect 168 604 171 612
rect 196 608 199 646
rect 253 538 256 653
rect 443 643 446 702
rect 443 640 462 643
rect 357 625 360 632
rect 459 633 462 640
rect 459 630 465 633
rect 357 622 456 625
rect 357 616 360 622
rect 329 613 360 616
rect 329 602 332 613
rect 341 605 381 608
rect 453 604 456 622
rect 270 599 332 602
rect 462 591 465 630
rect 459 588 465 591
rect 253 535 354 538
rect 157 527 332 530
rect -336 509 -262 512
rect -336 485 -333 509
rect -314 486 -273 489
rect -275 476 -259 479
rect -258 463 -255 474
rect -186 462 -183 475
rect -167 465 -164 526
rect -79 517 -67 520
rect -155 492 -115 495
rect -114 482 -110 492
rect 64 481 67 519
rect 225 498 228 505
rect 225 495 324 498
rect 225 489 228 495
rect 197 486 228 489
rect 197 475 200 486
rect 209 478 249 481
rect 321 477 324 495
rect 138 472 200 475
rect 329 469 332 527
rect 342 486 345 507
rect 351 496 354 535
rect 459 534 462 588
rect 480 581 483 721
rect 513 640 516 739
rect 555 648 558 686
rect 716 665 719 672
rect 820 671 823 728
rect 820 668 898 671
rect 716 662 815 665
rect 716 656 719 662
rect 688 653 719 656
rect 513 637 531 640
rect 688 642 691 653
rect 700 645 740 648
rect 812 644 815 662
rect 629 639 691 642
rect 480 578 686 581
rect 471 536 474 552
rect 374 531 462 534
rect 480 534 483 578
rect 494 561 521 564
rect 518 558 521 561
rect 518 557 534 558
rect 518 555 544 557
rect 531 554 669 555
rect 531 550 534 554
rect 541 552 669 554
rect 480 531 513 534
rect 480 522 483 531
rect 423 519 483 522
rect 329 466 341 469
rect -167 462 -151 465
rect 18 460 41 464
rect 22 389 26 460
rect 338 454 341 466
rect 250 451 348 454
rect 250 354 253 451
rect 332 413 335 431
rect 104 351 253 354
rect 260 410 335 413
rect 260 352 263 410
rect 345 406 348 451
rect 269 403 348 406
rect 269 363 272 403
rect 355 399 358 475
rect 279 396 358 399
rect 279 374 282 396
rect 363 391 366 488
rect 290 388 366 391
rect 290 384 293 388
rect -1271 303 -1014 306
rect -1271 251 -1268 303
rect -1301 248 -1259 251
rect -1311 239 -1285 242
rect -1261 238 -1245 241
rect -1245 225 -1240 236
rect -1172 224 -1169 237
rect -1153 227 -1150 288
rect -1065 279 -1053 282
rect -1141 254 -1101 257
rect -1100 244 -1096 254
rect -1153 224 -1137 227
rect -1017 205 -1014 303
rect -612 302 -355 305
rect -995 271 -921 274
rect -995 247 -992 271
rect -973 248 -932 251
rect -934 238 -918 241
rect -917 225 -914 236
rect -845 224 -842 237
rect -826 227 -823 288
rect -738 279 -726 282
rect -814 254 -774 257
rect -773 244 -769 254
rect -612 250 -609 302
rect -642 247 -600 250
rect -652 238 -626 241
rect -602 237 -586 240
rect -826 224 -810 227
rect -586 224 -581 235
rect -513 223 -510 236
rect -494 226 -491 287
rect -406 278 -394 281
rect -482 253 -442 256
rect -441 243 -437 253
rect -494 223 -478 226
rect -358 204 -355 302
rect 65 299 68 337
rect -336 270 -262 273
rect -336 246 -333 270
rect -314 247 -273 250
rect -275 237 -259 240
rect -258 224 -255 235
rect -186 223 -183 236
rect -167 226 -164 287
rect -79 278 -67 281
rect 19 278 42 282
rect -155 253 -115 256
rect -114 243 -110 253
rect -167 223 -151 226
rect 23 207 27 278
rect 104 221 107 351
rect 279 339 282 369
rect 113 336 282 339
rect 113 229 116 336
rect 226 316 229 323
rect 259 320 282 323
rect 259 316 262 320
rect 226 313 262 316
rect 279 316 282 320
rect 279 313 325 316
rect 226 307 229 313
rect 198 304 229 307
rect 198 293 201 304
rect 210 296 250 299
rect 139 290 201 293
rect 257 234 261 258
rect 270 233 274 305
rect 322 295 325 313
rect 113 226 237 229
rect 289 229 293 258
rect 104 218 230 221
rect 227 203 230 218
rect 234 216 237 226
rect 289 225 311 229
rect 330 226 333 388
rect 423 382 426 519
rect 497 488 500 517
rect 510 495 513 531
rect 510 492 526 495
rect 497 484 501 488
rect 499 471 512 474
rect 499 463 502 471
rect 459 460 502 463
rect 485 459 489 460
rect 494 400 498 441
rect 507 410 510 446
rect 656 439 660 485
rect 526 435 660 439
rect 666 448 669 552
rect 683 527 686 578
rect 683 524 857 527
rect 854 460 857 524
rect 854 454 857 455
rect 666 445 872 448
rect 526 400 530 435
rect 666 424 669 445
rect 854 432 857 433
rect 564 421 669 424
rect 494 398 499 400
rect 526 398 531 400
rect 494 394 531 398
rect 564 381 567 421
rect 656 403 695 406
rect 405 350 408 359
rect 656 359 659 403
rect 702 376 771 379
rect 768 365 771 376
rect 787 376 790 411
rect 824 400 826 404
rect 824 392 827 400
rect 824 389 835 392
rect 787 373 819 376
rect 832 365 835 389
rect 768 362 835 365
rect 372 347 408 350
rect 414 335 417 349
rect 555 352 558 358
rect 523 349 558 352
rect 689 341 692 351
rect 380 332 417 335
rect 689 338 706 341
rect 426 328 429 332
rect 570 328 573 336
rect 426 325 573 328
rect 426 318 429 325
rect 371 315 429 318
rect 705 320 708 329
rect 582 319 708 320
rect 562 317 708 319
rect 562 316 586 317
rect 462 301 465 315
rect 589 309 697 312
rect 589 301 592 309
rect 462 298 592 301
rect 839 291 842 413
rect 326 223 333 226
rect 337 288 842 291
rect 234 213 312 216
rect 227 200 280 203
rect 309 193 312 213
rect 326 201 329 223
rect 337 219 340 288
rect 854 273 857 427
rect 441 270 857 273
rect 388 230 391 268
rect 326 198 362 201
rect 309 190 354 193
rect -1271 116 -1014 119
rect -1271 64 -1268 116
rect -1301 61 -1259 64
rect -1311 52 -1285 55
rect -1261 51 -1245 54
rect -1245 38 -1240 49
rect -1172 37 -1169 50
rect -1153 40 -1150 101
rect -1065 92 -1053 95
rect -1141 67 -1101 70
rect -1100 57 -1096 67
rect -1153 37 -1137 40
rect -1017 18 -1014 116
rect -612 115 -355 118
rect 66 116 69 154
rect 227 133 230 140
rect 351 142 354 190
rect 359 151 362 198
rect 441 166 444 270
rect 869 261 872 445
rect 895 391 898 668
rect 901 330 925 334
rect 549 247 552 254
rect 655 258 872 261
rect 921 259 925 330
rect 549 244 648 247
rect 549 238 552 244
rect 521 235 552 238
rect 521 224 524 235
rect 533 227 573 230
rect 645 226 648 244
rect 462 221 524 224
rect 441 163 508 166
rect 359 148 363 151
rect 351 139 355 142
rect 360 140 363 148
rect 505 143 508 163
rect 655 159 658 258
rect 921 255 989 259
rect 673 243 812 247
rect 675 230 692 234
rect 1013 227 1016 265
rect 1174 244 1177 251
rect 1174 241 1273 244
rect 1174 235 1177 241
rect 1146 232 1177 235
rect 1146 221 1149 232
rect 1158 224 1198 227
rect 1270 223 1273 241
rect 1087 218 1149 221
rect 633 156 658 159
rect 227 130 326 133
rect 227 124 230 130
rect 199 121 230 124
rect -995 84 -921 87
rect -995 60 -992 84
rect -973 61 -932 64
rect -934 51 -918 54
rect -917 38 -914 49
rect -845 37 -842 50
rect -826 40 -823 101
rect -738 92 -726 95
rect -814 67 -774 70
rect -773 57 -769 67
rect -612 63 -609 115
rect -642 60 -600 63
rect -652 51 -626 54
rect -602 50 -586 53
rect -826 37 -810 40
rect -586 37 -581 48
rect -513 36 -510 49
rect -494 39 -491 100
rect -406 91 -394 94
rect -482 66 -442 69
rect -441 56 -437 66
rect -494 36 -478 39
rect -358 17 -355 115
rect 199 110 202 121
rect 211 113 251 116
rect 323 112 326 130
rect 140 107 202 110
rect 336 110 339 131
rect 352 129 355 139
rect 633 129 636 156
rect 352 127 360 129
rect 352 126 356 127
rect 487 121 494 124
rect 487 115 490 121
rect 455 112 490 115
rect 494 106 499 107
rect 455 103 499 106
rect 622 112 625 113
rect 590 109 625 112
rect -336 83 -262 86
rect -336 59 -333 83
rect -314 60 -273 63
rect -275 50 -259 53
rect -258 37 -255 48
rect -186 36 -183 49
rect -167 39 -164 100
rect 20 95 43 99
rect -79 91 -67 94
rect -155 66 -115 69
rect -114 56 -110 66
rect -167 36 -151 39
rect 24 24 28 95
rect 455 94 503 97
rect 599 99 624 102
rect 337 82 340 84
rect 309 79 340 82
rect 337 73 340 79
rect 512 80 515 84
rect 641 82 644 92
rect 665 82 668 174
rect 679 158 682 185
rect 817 169 820 200
rect 976 169 979 205
rect 817 166 979 169
rect 679 155 733 158
rect 730 114 733 155
rect 817 82 820 166
rect 831 98 835 127
rect 641 80 820 82
rect 512 79 820 80
rect 512 77 644 79
rect 512 73 515 77
rect 337 70 515 73
<< ntransistor >>
rect 660 1313 662 1333
rect 668 1313 670 1333
rect 725 1313 727 1333
rect 733 1313 735 1333
rect 802 1313 804 1333
rect 810 1313 812 1333
rect 867 1313 869 1333
rect 875 1313 877 1333
rect 942 1313 944 1333
rect 950 1313 952 1333
rect 1007 1313 1009 1333
rect 1015 1313 1017 1333
rect 1087 1313 1089 1333
rect 1095 1313 1097 1333
rect 1152 1313 1154 1333
rect 1160 1313 1162 1333
rect 1232 1313 1234 1333
rect 1240 1313 1242 1333
rect 1297 1313 1299 1333
rect 1305 1313 1307 1333
rect 1377 1313 1379 1333
rect 1385 1313 1387 1333
rect 1442 1313 1444 1333
rect 1450 1313 1452 1333
rect 678 1207 680 1227
rect 686 1207 688 1227
rect 725 1207 727 1227
rect 733 1207 735 1227
rect 820 1207 822 1227
rect 828 1207 830 1227
rect 867 1207 869 1227
rect 875 1207 877 1227
rect 960 1207 962 1227
rect 968 1207 970 1227
rect 1007 1207 1009 1227
rect 1015 1207 1017 1227
rect 1105 1207 1107 1227
rect 1113 1207 1115 1227
rect 1152 1207 1154 1227
rect 1160 1207 1162 1227
rect 1250 1207 1252 1227
rect 1258 1207 1260 1227
rect 1297 1207 1299 1227
rect 1305 1207 1307 1227
rect 1395 1207 1397 1227
rect 1403 1207 1405 1227
rect 1442 1207 1444 1227
rect 1450 1207 1452 1227
rect -432 1127 -412 1129
rect 739 1131 749 1133
rect 881 1131 891 1133
rect 1021 1131 1031 1133
rect 1166 1131 1176 1133
rect 1311 1131 1321 1133
rect 1456 1131 1466 1133
rect -105 1127 -85 1129
rect -432 1119 -412 1121
rect -105 1119 -85 1121
rect -538 1109 -518 1111
rect -211 1109 -191 1111
rect -538 1101 -518 1103
rect -211 1101 -191 1103
rect -538 1062 -518 1064
rect 739 1081 749 1083
rect 881 1081 891 1083
rect 1021 1081 1031 1083
rect 1166 1081 1176 1083
rect 1311 1081 1321 1083
rect 1456 1081 1466 1083
rect -432 1062 -412 1064
rect -538 1054 -518 1056
rect -665 1040 -663 1050
rect -614 1040 -612 1050
rect -432 1054 -412 1056
rect -211 1062 -191 1064
rect -105 1062 -85 1064
rect -211 1054 -191 1056
rect -337 1040 -335 1050
rect -287 1040 -285 1050
rect -105 1054 -85 1056
rect 452 1025 472 1027
rect 452 1017 472 1019
rect 361 991 381 993
rect 548 991 568 993
rect 361 983 381 985
rect 660 986 662 1006
rect 668 986 670 1006
rect 725 986 727 1006
rect 733 986 735 1006
rect 802 986 804 1006
rect 810 986 812 1006
rect 867 986 869 1006
rect 875 986 877 1006
rect 942 986 944 1006
rect 950 986 952 1006
rect 1007 986 1009 1006
rect 1015 986 1017 1006
rect 1087 986 1089 1006
rect 1095 986 1097 1006
rect 1152 986 1154 1006
rect 1160 986 1162 1006
rect 1232 986 1234 1006
rect 1240 986 1242 1006
rect 1297 986 1299 1006
rect 1305 986 1307 1006
rect 1377 986 1379 1006
rect 1385 986 1387 1006
rect 1442 986 1444 1006
rect 1450 986 1452 1006
rect 548 983 568 985
rect -1092 967 -1072 969
rect -765 967 -745 969
rect -1092 959 -1072 961
rect -433 963 -413 965
rect -765 959 -745 961
rect -1198 949 -1178 951
rect 452 969 472 971
rect -106 963 -86 965
rect -433 955 -413 957
rect -871 949 -851 951
rect -1198 941 -1178 943
rect 452 961 472 963
rect -106 955 -86 957
rect -539 945 -519 947
rect -871 941 -851 943
rect -212 945 -192 947
rect -539 937 -519 939
rect -212 937 -192 939
rect 201 937 221 939
rect 201 929 221 931
rect -1198 902 -1178 904
rect -1092 902 -1072 904
rect -1198 894 -1178 896
rect -1325 880 -1323 890
rect -1274 880 -1272 890
rect -1092 894 -1072 896
rect -871 902 -851 904
rect -765 902 -745 904
rect -871 894 -851 896
rect -997 880 -995 890
rect -947 880 -945 890
rect -765 894 -745 896
rect -539 898 -519 900
rect -433 898 -413 900
rect -539 890 -519 892
rect -666 876 -664 886
rect -615 876 -613 886
rect -433 890 -413 892
rect -212 898 -192 900
rect 110 903 130 905
rect -106 898 -86 900
rect -212 890 -192 892
rect -338 876 -336 886
rect -288 876 -286 886
rect 297 903 317 905
rect 110 895 130 897
rect -106 890 -86 892
rect 297 895 317 897
rect 401 884 421 886
rect 201 881 221 883
rect 401 876 421 878
rect 538 883 548 885
rect 201 873 221 875
rect 446 866 448 876
rect 538 875 548 877
rect 678 880 680 900
rect 686 880 688 900
rect 725 880 727 900
rect 733 880 735 900
rect 820 880 822 900
rect 828 880 830 900
rect 867 880 869 900
rect 875 880 877 900
rect 960 880 962 900
rect 968 880 970 900
rect 1007 880 1009 900
rect 1015 880 1017 900
rect 1105 880 1107 900
rect 1113 880 1115 900
rect 1152 880 1154 900
rect 1160 880 1162 900
rect 1250 880 1252 900
rect 1258 880 1260 900
rect 1297 880 1299 900
rect 1305 880 1307 900
rect 1395 880 1397 900
rect 1403 880 1405 900
rect 1442 880 1444 900
rect 1450 880 1452 900
rect 574 866 576 876
rect 92 823 112 825
rect 92 815 112 817
rect 137 805 139 815
rect 324 798 344 800
rect 324 790 344 792
rect 487 801 497 803
rect 739 804 749 806
rect 881 804 891 806
rect 1021 804 1031 806
rect 1166 804 1176 806
rect 1311 804 1321 806
rect 1456 804 1466 806
rect 487 793 497 795
rect 369 780 371 790
rect 487 785 497 787
rect 522 773 524 783
rect 200 757 220 759
rect 739 753 749 755
rect 881 753 891 755
rect 1021 753 1031 755
rect 1166 753 1176 755
rect 1311 753 1321 755
rect 1456 753 1466 755
rect 200 749 220 751
rect -1092 728 -1072 730
rect -765 728 -745 730
rect -1092 720 -1072 722
rect -433 727 -413 729
rect -765 720 -745 722
rect -1198 710 -1178 712
rect -106 727 -86 729
rect -433 719 -413 721
rect -871 710 -851 712
rect -1198 702 -1178 704
rect 109 723 129 725
rect -106 719 -86 721
rect -539 709 -519 711
rect -871 702 -851 704
rect 296 723 316 725
rect 109 715 129 717
rect -212 709 -192 711
rect 296 715 316 717
rect 406 716 436 718
rect -539 701 -519 703
rect -212 701 -192 703
rect 406 708 436 710
rect 200 701 220 703
rect 406 700 436 702
rect 200 693 220 695
rect 461 687 463 697
rect -1198 663 -1178 665
rect -1092 663 -1072 665
rect -1198 655 -1178 657
rect -1325 641 -1323 651
rect -1274 641 -1272 651
rect -1092 655 -1072 657
rect -871 663 -851 665
rect -765 663 -745 665
rect -871 655 -851 657
rect -997 641 -995 651
rect -947 641 -945 651
rect -765 655 -745 657
rect -539 662 -519 664
rect -433 662 -413 664
rect -539 654 -519 656
rect -666 640 -664 650
rect -615 640 -613 650
rect -433 654 -413 656
rect -212 662 -192 664
rect -106 662 -86 664
rect -212 654 -192 656
rect -338 640 -336 650
rect -288 640 -286 650
rect -106 654 -86 656
rect 691 670 711 672
rect 691 662 711 664
rect 91 643 111 645
rect 91 635 111 637
rect 136 625 138 635
rect 600 636 620 638
rect 332 630 352 632
rect 787 636 807 638
rect 600 628 620 630
rect 332 622 352 624
rect 787 628 807 630
rect 691 614 711 616
rect 691 606 711 608
rect 241 596 261 598
rect 428 596 448 598
rect 241 588 261 590
rect 428 588 448 590
rect 332 574 352 576
rect 332 566 352 568
rect 581 532 601 534
rect 581 524 601 526
rect -1092 514 -1072 516
rect -765 514 -745 516
rect -1092 506 -1072 508
rect -433 513 -413 515
rect -765 506 -745 508
rect -1198 496 -1178 498
rect -106 513 -86 515
rect 626 514 628 524
rect -433 505 -413 507
rect -871 496 -851 498
rect -1198 488 -1178 490
rect -106 505 -86 507
rect -539 495 -519 497
rect -871 488 -851 490
rect 200 503 220 505
rect -212 495 -192 497
rect -539 487 -519 489
rect 200 495 220 497
rect -212 487 -192 489
rect 411 481 451 483
rect -1198 449 -1178 451
rect -1092 449 -1072 451
rect -1198 441 -1178 443
rect -1325 427 -1323 437
rect -1274 427 -1272 437
rect -1092 441 -1072 443
rect -871 449 -851 451
rect -765 449 -745 451
rect -871 441 -851 443
rect -997 427 -995 437
rect -947 427 -945 437
rect -765 441 -745 443
rect -539 448 -519 450
rect 109 469 129 471
rect 580 479 610 481
rect 411 473 451 475
rect 296 469 316 471
rect 109 461 129 463
rect 411 465 451 467
rect 296 461 316 463
rect 787 495 797 497
rect 787 487 797 489
rect 787 479 797 481
rect 580 471 610 473
rect 580 463 610 465
rect 411 457 451 459
rect -433 448 -413 450
rect -539 440 -519 442
rect -666 426 -664 436
rect -615 426 -613 436
rect -433 440 -413 442
rect -212 448 -192 450
rect -106 448 -86 450
rect -212 440 -192 442
rect -338 426 -336 436
rect -288 426 -286 436
rect 476 449 478 459
rect 787 471 797 473
rect 823 461 825 471
rect 635 450 637 460
rect 200 447 220 449
rect -106 440 -86 442
rect 200 439 220 441
rect 758 411 778 413
rect 758 403 778 405
rect 91 389 111 391
rect 91 381 111 383
rect 803 393 805 403
rect 136 371 138 381
rect 339 368 364 370
rect 475 370 515 372
rect 339 360 364 362
rect 339 352 364 354
rect 621 367 651 369
rect 475 362 515 364
rect 475 354 515 356
rect 339 344 364 346
rect 339 336 364 338
rect 390 337 392 347
rect 621 359 651 361
rect 621 351 651 353
rect 475 346 515 348
rect 540 338 542 348
rect 676 338 678 348
rect 847 347 857 349
rect 847 339 857 341
rect 847 331 857 333
rect 201 321 221 323
rect 847 323 857 325
rect 201 313 221 315
rect 881 317 883 327
rect 847 315 857 317
rect 110 287 130 289
rect -1092 275 -1072 277
rect -765 275 -745 277
rect -1092 267 -1072 269
rect -433 274 -413 276
rect -765 267 -745 269
rect -1198 257 -1178 259
rect 297 287 317 289
rect 110 279 130 281
rect -106 274 -86 276
rect 297 279 317 281
rect -433 266 -413 268
rect -871 257 -851 259
rect -1198 249 -1178 251
rect -106 266 -86 268
rect -539 256 -519 258
rect -871 249 -851 251
rect 201 265 221 267
rect -212 256 -192 258
rect 201 257 221 259
rect -539 248 -519 250
rect 524 252 544 254
rect -212 248 -192 250
rect 1149 249 1169 251
rect 524 244 544 246
rect 1149 241 1169 243
rect -1198 210 -1178 212
rect -1092 210 -1072 212
rect -1198 202 -1178 204
rect -1325 188 -1323 198
rect -1274 188 -1272 198
rect -1092 202 -1072 204
rect -871 210 -851 212
rect -765 210 -745 212
rect -871 202 -851 204
rect -997 188 -995 198
rect -947 188 -945 198
rect -765 202 -745 204
rect -539 209 -519 211
rect -433 209 -413 211
rect -539 201 -519 203
rect -666 187 -664 197
rect -615 187 -613 197
rect -433 201 -413 203
rect -212 209 -192 211
rect 433 218 453 220
rect -106 209 -86 211
rect -212 201 -192 203
rect -338 187 -336 197
rect -288 187 -286 197
rect 92 207 112 209
rect -106 201 -86 203
rect 92 199 112 201
rect 620 218 640 220
rect 433 210 453 212
rect 620 210 640 212
rect 137 189 139 199
rect 738 199 768 201
rect 524 196 544 198
rect 885 211 905 213
rect 885 203 905 205
rect 1058 215 1078 217
rect 1245 215 1265 217
rect 1058 207 1078 209
rect 738 191 768 193
rect 524 188 544 190
rect 738 183 768 185
rect 930 193 932 203
rect 1245 207 1265 209
rect 1149 193 1169 195
rect 1149 185 1169 187
rect 793 170 795 180
rect 202 138 222 140
rect 202 130 222 132
rect 413 128 443 130
rect 413 120 443 122
rect 557 130 582 132
rect 557 122 582 124
rect 413 112 443 114
rect 111 104 131 106
rect 298 104 318 106
rect 111 96 131 98
rect -1092 88 -1072 90
rect -765 88 -745 90
rect -1092 80 -1072 82
rect -433 87 -413 89
rect -765 80 -745 82
rect -1198 70 -1178 72
rect 413 104 443 106
rect 298 96 318 98
rect 557 114 582 116
rect 685 122 725 124
rect 996 126 1006 128
rect 996 118 1006 120
rect 685 114 725 116
rect 557 106 582 108
rect 413 96 443 98
rect -106 87 -86 89
rect -433 79 -413 81
rect -871 70 -851 72
rect -1198 62 -1178 64
rect 475 90 477 100
rect 557 98 582 100
rect 608 99 610 109
rect 685 106 725 108
rect 996 110 1006 112
rect 996 102 1006 104
rect 685 98 725 100
rect 750 90 752 100
rect 996 94 1006 96
rect 413 88 443 90
rect 202 82 222 84
rect 1039 88 1041 98
rect 996 86 1006 88
rect -106 79 -86 81
rect -539 69 -519 71
rect -871 62 -851 64
rect 202 74 222 76
rect -212 69 -192 71
rect -539 61 -519 63
rect -212 61 -192 63
rect -1198 23 -1178 25
rect -1092 23 -1072 25
rect -1198 15 -1178 17
rect -1325 1 -1323 11
rect -1274 1 -1272 11
rect -1092 15 -1072 17
rect -871 23 -851 25
rect -765 23 -745 25
rect -871 15 -851 17
rect -997 1 -995 11
rect -947 1 -945 11
rect -765 15 -745 17
rect -539 22 -519 24
rect -433 22 -413 24
rect -539 14 -519 16
rect -666 0 -664 10
rect -615 0 -613 10
rect -433 14 -413 16
rect -212 22 -192 24
rect -106 22 -86 24
rect 93 24 113 26
rect -212 14 -192 16
rect -338 0 -336 10
rect -288 0 -286 10
rect -106 14 -86 16
rect 93 16 113 18
rect 138 6 140 16
<< ptransistor >>
rect 660 1277 662 1297
rect 668 1277 670 1297
rect 725 1277 727 1297
rect 733 1277 735 1297
rect 802 1277 804 1297
rect 810 1277 812 1297
rect 867 1277 869 1297
rect 875 1277 877 1297
rect 942 1277 944 1297
rect 950 1277 952 1297
rect 1007 1277 1009 1297
rect 1015 1277 1017 1297
rect 1087 1277 1089 1297
rect 1095 1277 1097 1297
rect 1152 1277 1154 1297
rect 1160 1277 1162 1297
rect 1232 1277 1234 1297
rect 1240 1277 1242 1297
rect 1297 1277 1299 1297
rect 1305 1277 1307 1297
rect 1377 1277 1379 1297
rect 1385 1277 1387 1297
rect 1442 1277 1444 1297
rect 1450 1277 1452 1297
rect 678 1171 680 1191
rect 686 1171 688 1191
rect 725 1171 727 1191
rect 733 1171 735 1191
rect 820 1171 822 1191
rect 828 1171 830 1191
rect 867 1171 869 1191
rect 875 1171 877 1191
rect 960 1171 962 1191
rect 968 1171 970 1191
rect 1007 1171 1009 1191
rect 1015 1171 1017 1191
rect 1105 1171 1107 1191
rect 1113 1171 1115 1191
rect 1152 1171 1154 1191
rect 1160 1171 1162 1191
rect 1250 1171 1252 1191
rect 1258 1171 1260 1191
rect 1297 1171 1299 1191
rect 1305 1171 1307 1191
rect 1395 1171 1397 1191
rect 1403 1171 1405 1191
rect 1442 1171 1444 1191
rect 1450 1171 1452 1191
rect -468 1127 -448 1129
rect 705 1131 725 1133
rect 847 1131 867 1133
rect 987 1131 1007 1133
rect 1132 1131 1152 1133
rect 1277 1131 1297 1133
rect 1422 1131 1442 1133
rect -141 1127 -121 1129
rect -468 1119 -448 1121
rect -141 1119 -121 1121
rect -574 1109 -554 1111
rect -247 1109 -227 1111
rect -574 1101 -554 1103
rect -247 1101 -227 1103
rect -665 1064 -663 1084
rect -614 1064 -612 1084
rect -574 1062 -554 1064
rect -337 1064 -335 1084
rect -287 1064 -285 1084
rect 705 1081 725 1083
rect 847 1081 867 1083
rect 987 1081 1007 1083
rect 1132 1081 1152 1083
rect 1277 1081 1297 1083
rect 1422 1081 1442 1083
rect -468 1062 -448 1064
rect -574 1054 -554 1056
rect -468 1054 -448 1056
rect -247 1062 -227 1064
rect -141 1062 -121 1064
rect -247 1054 -227 1056
rect -141 1054 -121 1056
rect 416 1025 436 1027
rect 416 1017 436 1019
rect 325 991 345 993
rect 512 991 532 993
rect 325 983 345 985
rect 512 983 532 985
rect -1128 967 -1108 969
rect -801 967 -781 969
rect -1128 959 -1108 961
rect -469 963 -449 965
rect -801 959 -781 961
rect -1234 949 -1214 951
rect 416 969 436 971
rect -142 963 -122 965
rect -469 955 -449 957
rect -907 949 -887 951
rect -1234 941 -1214 943
rect 416 961 436 963
rect -142 955 -122 957
rect -575 945 -555 947
rect -907 941 -887 943
rect 660 950 662 970
rect 668 950 670 970
rect 725 950 727 970
rect 733 950 735 970
rect 802 950 804 970
rect 810 950 812 970
rect 867 950 869 970
rect 875 950 877 970
rect 942 950 944 970
rect 950 950 952 970
rect 1007 950 1009 970
rect 1015 950 1017 970
rect 1087 950 1089 970
rect 1095 950 1097 970
rect 1152 950 1154 970
rect 1160 950 1162 970
rect 1232 950 1234 970
rect 1240 950 1242 970
rect 1297 950 1299 970
rect 1305 950 1307 970
rect 1377 950 1379 970
rect 1385 950 1387 970
rect 1442 950 1444 970
rect 1450 950 1452 970
rect -248 945 -228 947
rect -575 937 -555 939
rect -248 937 -228 939
rect 165 937 185 939
rect 165 929 185 931
rect -1325 904 -1323 924
rect -1274 904 -1272 924
rect -1234 902 -1214 904
rect -997 904 -995 924
rect -947 904 -945 924
rect -1128 902 -1108 904
rect -1234 894 -1214 896
rect -1128 894 -1108 896
rect -907 902 -887 904
rect -801 902 -781 904
rect -907 894 -887 896
rect -666 900 -664 920
rect -615 900 -613 920
rect -801 894 -781 896
rect -575 898 -555 900
rect -338 900 -336 920
rect -288 900 -286 920
rect -469 898 -449 900
rect -575 890 -555 892
rect -469 890 -449 892
rect -248 898 -228 900
rect 74 903 94 905
rect -142 898 -122 900
rect -248 890 -228 892
rect 261 903 281 905
rect 74 895 94 897
rect -142 890 -122 892
rect 261 895 281 897
rect 446 892 448 912
rect 574 892 576 912
rect 368 884 388 886
rect 165 881 185 883
rect 368 876 388 878
rect 486 883 526 885
rect 165 873 185 875
rect 486 875 526 877
rect 137 831 139 851
rect 678 844 680 864
rect 686 844 688 864
rect 725 844 727 864
rect 733 844 735 864
rect 820 844 822 864
rect 828 844 830 864
rect 867 844 869 864
rect 875 844 877 864
rect 960 844 962 864
rect 968 844 970 864
rect 1007 844 1009 864
rect 1015 844 1017 864
rect 1105 844 1107 864
rect 1113 844 1115 864
rect 1152 844 1154 864
rect 1160 844 1162 864
rect 1250 844 1252 864
rect 1258 844 1260 864
rect 1297 844 1299 864
rect 1305 844 1307 864
rect 1395 844 1397 864
rect 1403 844 1405 864
rect 1442 844 1444 864
rect 1450 844 1452 864
rect 59 823 79 825
rect 59 815 79 817
rect 369 806 371 826
rect 291 798 311 800
rect 291 790 311 792
rect 415 801 475 803
rect 522 799 524 819
rect 705 804 725 806
rect 847 804 867 806
rect 987 804 1007 806
rect 1132 804 1152 806
rect 1277 804 1297 806
rect 1422 804 1442 806
rect 415 793 475 795
rect 415 785 475 787
rect 164 757 184 759
rect 705 753 725 755
rect 847 753 867 755
rect 987 753 1007 755
rect 1132 753 1152 755
rect 1277 753 1297 755
rect 1422 753 1442 755
rect 164 749 184 751
rect -1128 728 -1108 730
rect -801 728 -781 730
rect -1128 720 -1108 722
rect -469 727 -449 729
rect -801 720 -781 722
rect -1234 710 -1214 712
rect -142 727 -122 729
rect -469 719 -449 721
rect -907 710 -887 712
rect -1234 702 -1214 704
rect 73 723 93 725
rect -142 719 -122 721
rect -575 709 -555 711
rect -907 702 -887 704
rect 260 723 280 725
rect 73 715 93 717
rect -248 709 -228 711
rect 260 715 280 717
rect 374 716 394 718
rect -575 701 -555 703
rect -248 701 -228 703
rect 461 713 463 733
rect 374 708 394 710
rect 164 701 184 703
rect 374 700 394 702
rect 164 693 184 695
rect -1325 665 -1323 685
rect -1274 665 -1272 685
rect -1234 663 -1214 665
rect -997 665 -995 685
rect -947 665 -945 685
rect -1128 663 -1108 665
rect -1234 655 -1214 657
rect -1128 655 -1108 657
rect -907 663 -887 665
rect -801 663 -781 665
rect -666 664 -664 684
rect -615 664 -613 684
rect -907 655 -887 657
rect -801 655 -781 657
rect -575 662 -555 664
rect -338 664 -336 684
rect -288 664 -286 684
rect -469 662 -449 664
rect -575 654 -555 656
rect -469 654 -449 656
rect -248 662 -228 664
rect -142 662 -122 664
rect -248 654 -228 656
rect -142 654 -122 656
rect 136 651 138 671
rect 655 670 675 672
rect 655 662 675 664
rect 58 643 78 645
rect 58 635 78 637
rect 564 636 584 638
rect 296 630 316 632
rect 751 636 771 638
rect 564 628 584 630
rect 296 622 316 624
rect 751 628 771 630
rect 655 614 675 616
rect 655 606 675 608
rect 205 596 225 598
rect 392 596 412 598
rect 205 588 225 590
rect 392 588 412 590
rect 296 574 316 576
rect 296 566 316 568
rect 626 540 628 560
rect 548 532 568 534
rect 548 524 568 526
rect -1128 514 -1108 516
rect -801 514 -781 516
rect -1128 506 -1108 508
rect -469 513 -449 515
rect -801 506 -781 508
rect -1234 496 -1214 498
rect -142 513 -122 515
rect -469 505 -449 507
rect -907 496 -887 498
rect -1234 488 -1214 490
rect -142 505 -122 507
rect -575 495 -555 497
rect -907 488 -887 490
rect 164 503 184 505
rect -248 495 -228 497
rect -575 487 -555 489
rect 164 495 184 497
rect -248 487 -228 489
rect 379 481 399 483
rect -1325 451 -1323 471
rect -1274 451 -1272 471
rect -1234 449 -1214 451
rect -997 451 -995 471
rect -947 451 -945 471
rect -1128 449 -1108 451
rect -1234 441 -1214 443
rect -1128 441 -1108 443
rect -907 449 -887 451
rect -801 449 -781 451
rect -666 450 -664 470
rect -615 450 -613 470
rect -907 441 -887 443
rect -801 441 -781 443
rect -575 448 -555 450
rect -338 450 -336 470
rect -288 450 -286 470
rect 73 469 93 471
rect 476 475 478 495
rect 548 479 568 481
rect 379 473 399 475
rect 260 469 280 471
rect 73 461 93 463
rect 379 465 399 467
rect 260 461 280 463
rect 635 476 637 496
rect 695 495 775 497
rect 695 487 775 489
rect 823 487 825 507
rect 695 479 775 481
rect 548 471 568 473
rect 548 463 568 465
rect 379 457 399 459
rect -469 448 -449 450
rect -575 440 -555 442
rect -469 440 -449 442
rect -248 448 -228 450
rect -142 448 -122 450
rect -248 440 -228 442
rect 695 471 775 473
rect 164 447 184 449
rect -142 440 -122 442
rect 164 439 184 441
rect 803 419 805 439
rect 136 397 138 417
rect 725 411 745 413
rect 725 403 745 405
rect 58 389 78 391
rect 58 381 78 383
rect 307 368 327 370
rect 390 363 392 383
rect 443 370 463 372
rect 307 360 327 362
rect 307 352 327 354
rect 540 364 542 384
rect 589 367 609 369
rect 443 362 463 364
rect 443 354 463 356
rect 307 344 327 346
rect 307 336 327 338
rect 676 364 678 384
rect 589 359 609 361
rect 589 351 609 353
rect 443 346 463 348
rect 735 347 835 349
rect 881 343 883 363
rect 735 339 835 341
rect 735 331 835 333
rect 165 321 185 323
rect 735 323 835 325
rect 165 313 185 315
rect 735 315 835 317
rect 74 287 94 289
rect -1128 275 -1108 277
rect -801 275 -781 277
rect -1128 267 -1108 269
rect -469 274 -449 276
rect -801 267 -781 269
rect -1234 257 -1214 259
rect 261 287 281 289
rect 74 279 94 281
rect -142 274 -122 276
rect 261 279 281 281
rect -469 266 -449 268
rect -907 257 -887 259
rect -1234 249 -1214 251
rect -142 266 -122 268
rect -575 256 -555 258
rect -907 249 -887 251
rect 165 265 185 267
rect -248 256 -228 258
rect 165 257 185 259
rect -575 248 -555 250
rect 488 252 508 254
rect -248 248 -228 250
rect 1113 249 1133 251
rect 488 244 508 246
rect 1113 241 1133 243
rect -1325 212 -1323 232
rect -1274 212 -1272 232
rect -1234 210 -1214 212
rect -997 212 -995 232
rect -947 212 -945 232
rect -1128 210 -1108 212
rect -1234 202 -1214 204
rect -1128 202 -1108 204
rect -907 210 -887 212
rect -801 210 -781 212
rect -666 211 -664 231
rect -615 211 -613 231
rect -907 202 -887 204
rect -801 202 -781 204
rect -575 209 -555 211
rect -338 211 -336 231
rect -288 211 -286 231
rect -469 209 -449 211
rect -575 201 -555 203
rect -469 201 -449 203
rect -248 209 -228 211
rect 137 215 139 235
rect 397 218 417 220
rect -142 209 -122 211
rect -248 201 -228 203
rect 59 207 79 209
rect -142 201 -122 203
rect 59 199 79 201
rect 584 218 604 220
rect 930 219 932 239
rect 397 210 417 212
rect 584 210 604 212
rect 706 199 726 201
rect 488 196 508 198
rect 793 196 795 216
rect 852 211 872 213
rect 852 203 872 205
rect 1022 215 1042 217
rect 1209 215 1229 217
rect 1022 207 1042 209
rect 706 191 726 193
rect 488 188 508 190
rect 706 183 726 185
rect 1209 207 1229 209
rect 1113 193 1133 195
rect 1113 185 1133 187
rect 166 138 186 140
rect 166 130 186 132
rect 389 128 399 130
rect 389 120 399 122
rect 475 116 477 136
rect 525 130 545 132
rect 608 125 610 145
rect 525 122 545 124
rect 389 112 399 114
rect 75 104 95 106
rect 262 104 282 106
rect 75 96 95 98
rect -1128 88 -1108 90
rect -801 88 -781 90
rect -1128 80 -1108 82
rect -469 87 -449 89
rect -801 80 -781 82
rect -1234 70 -1214 72
rect 389 104 399 106
rect 262 96 282 98
rect 525 114 545 116
rect 653 122 673 124
rect 750 116 752 136
rect 864 126 984 128
rect 864 118 984 120
rect 653 114 673 116
rect 525 106 545 108
rect 389 96 399 98
rect -142 87 -122 89
rect -469 79 -449 81
rect -907 70 -887 72
rect -1234 62 -1214 64
rect 525 98 545 100
rect 653 106 673 108
rect 1039 114 1041 134
rect 864 110 984 112
rect 864 102 984 104
rect 653 98 673 100
rect 864 94 984 96
rect 389 88 399 90
rect 166 82 186 84
rect 864 86 984 88
rect -142 79 -122 81
rect -575 69 -555 71
rect -907 62 -887 64
rect 166 74 186 76
rect -248 69 -228 71
rect -575 61 -555 63
rect -248 61 -228 63
rect -1325 25 -1323 45
rect -1274 25 -1272 45
rect -1234 23 -1214 25
rect -997 25 -995 45
rect -947 25 -945 45
rect -1128 23 -1108 25
rect -1234 15 -1214 17
rect -1128 15 -1108 17
rect -907 23 -887 25
rect -801 23 -781 25
rect -666 24 -664 44
rect -615 24 -613 44
rect -907 15 -887 17
rect -801 15 -781 17
rect -575 22 -555 24
rect -338 24 -336 44
rect -288 24 -286 44
rect 138 32 140 52
rect -469 22 -449 24
rect -575 14 -555 16
rect -469 14 -449 16
rect -248 22 -228 24
rect -142 22 -122 24
rect 60 24 80 26
rect -248 14 -228 16
rect -142 14 -122 16
rect 60 16 80 18
<< polycontact >>
rect 659 1261 663 1265
rect 667 1261 671 1265
rect 724 1261 728 1265
rect 732 1261 736 1265
rect 801 1261 805 1265
rect 809 1261 813 1265
rect 866 1261 870 1265
rect 874 1261 878 1265
rect 941 1261 945 1265
rect 949 1261 953 1265
rect 1006 1261 1010 1265
rect 1014 1261 1018 1265
rect 1086 1261 1090 1265
rect 1094 1261 1098 1265
rect 1151 1261 1155 1265
rect 1159 1261 1163 1265
rect 1231 1261 1235 1265
rect 1239 1261 1243 1265
rect 1296 1261 1300 1265
rect 1304 1261 1308 1265
rect 1376 1261 1380 1265
rect 1384 1261 1388 1265
rect 1441 1261 1445 1265
rect 1449 1261 1453 1265
rect 677 1155 681 1159
rect 685 1155 689 1159
rect 724 1155 728 1159
rect 732 1155 736 1159
rect 819 1155 823 1159
rect 827 1155 831 1159
rect 866 1155 870 1159
rect 874 1155 878 1159
rect 959 1155 963 1159
rect 967 1155 971 1159
rect 1006 1155 1010 1159
rect 1014 1155 1018 1159
rect 1104 1155 1108 1159
rect 1112 1155 1116 1159
rect 1151 1155 1155 1159
rect 1159 1155 1163 1159
rect 1249 1155 1253 1159
rect 1257 1155 1261 1159
rect 1296 1155 1300 1159
rect 1304 1155 1308 1159
rect 1394 1155 1398 1159
rect 1402 1155 1406 1159
rect 1441 1155 1445 1159
rect 1449 1155 1453 1159
rect -484 1126 -480 1130
rect -484 1118 -480 1122
rect -157 1126 -153 1130
rect -590 1108 -586 1112
rect -157 1118 -153 1122
rect 732 1127 736 1131
rect 874 1127 878 1131
rect 1014 1127 1018 1131
rect 1159 1127 1163 1131
rect 1304 1127 1308 1131
rect 1449 1127 1453 1131
rect -590 1100 -586 1104
rect -263 1108 -259 1112
rect -263 1100 -259 1104
rect -669 1053 -665 1057
rect -618 1053 -614 1057
rect -590 1061 -586 1065
rect -590 1053 -586 1057
rect -484 1061 -480 1065
rect 732 1077 736 1081
rect 874 1077 878 1081
rect 1014 1077 1018 1081
rect 1159 1077 1163 1081
rect 1304 1077 1308 1081
rect 1449 1077 1453 1081
rect -484 1053 -480 1057
rect -341 1053 -337 1057
rect -291 1053 -287 1057
rect -263 1061 -259 1065
rect -263 1053 -259 1057
rect -157 1061 -153 1065
rect -157 1053 -153 1057
rect 400 1024 404 1028
rect 400 1016 404 1020
rect 309 990 313 994
rect 309 982 313 986
rect 496 990 500 994
rect 496 982 500 986
rect -1144 966 -1140 970
rect -1144 958 -1140 962
rect -817 966 -813 970
rect -1250 948 -1246 952
rect -817 958 -813 962
rect -485 962 -481 966
rect -1250 940 -1246 944
rect -923 948 -919 952
rect -485 954 -481 958
rect -158 962 -154 966
rect 400 968 404 972
rect -923 940 -919 944
rect -591 944 -587 948
rect -158 954 -154 958
rect 400 960 404 964
rect -591 936 -587 940
rect -264 944 -260 948
rect -264 936 -260 940
rect 149 936 153 940
rect 149 928 153 932
rect 659 934 663 938
rect 667 934 671 938
rect 724 934 728 938
rect 732 934 736 938
rect 801 934 805 938
rect 809 934 813 938
rect 866 934 870 938
rect 874 934 878 938
rect 941 934 945 938
rect 949 934 953 938
rect 1006 934 1010 938
rect 1014 934 1018 938
rect 1086 934 1090 938
rect 1094 934 1098 938
rect 1151 934 1155 938
rect 1159 934 1163 938
rect 1231 934 1235 938
rect 1239 934 1243 938
rect 1296 934 1300 938
rect 1304 934 1308 938
rect 1376 934 1380 938
rect 1384 934 1388 938
rect 1441 934 1445 938
rect 1449 934 1453 938
rect -1329 893 -1325 897
rect -1278 893 -1274 897
rect -1250 901 -1246 905
rect -1250 893 -1246 897
rect -1144 901 -1140 905
rect -1144 893 -1140 897
rect -1001 893 -997 897
rect -951 893 -947 897
rect -923 901 -919 905
rect -923 893 -919 897
rect -817 901 -813 905
rect -817 893 -813 897
rect -670 889 -666 893
rect -619 889 -615 893
rect -591 897 -587 901
rect -591 889 -587 893
rect -485 897 -481 901
rect -485 889 -481 893
rect -342 889 -338 893
rect -292 889 -288 893
rect -264 897 -260 901
rect -264 889 -260 893
rect -158 897 -154 901
rect 58 902 62 906
rect -158 889 -154 893
rect 58 894 62 898
rect 245 902 249 906
rect 245 894 249 898
rect 149 880 153 884
rect 355 883 359 887
rect 149 872 153 876
rect 355 875 359 879
rect 442 879 446 883
rect 473 882 477 886
rect 473 874 477 878
rect 570 879 574 883
rect 46 822 50 826
rect 46 814 50 818
rect 133 818 137 822
rect 677 828 681 832
rect 685 828 689 832
rect 724 828 728 832
rect 732 828 736 832
rect 819 828 823 832
rect 827 828 831 832
rect 866 828 870 832
rect 874 828 878 832
rect 959 828 963 832
rect 967 828 971 832
rect 1006 828 1010 832
rect 1014 828 1018 832
rect 1104 828 1108 832
rect 1112 828 1116 832
rect 1151 828 1155 832
rect 1159 828 1163 832
rect 1249 828 1253 832
rect 1257 828 1261 832
rect 1296 828 1300 832
rect 1304 828 1308 832
rect 1394 828 1398 832
rect 1402 828 1406 832
rect 1441 828 1445 832
rect 1449 828 1453 832
rect 278 797 282 801
rect 278 789 282 793
rect 365 793 369 797
rect 402 800 406 804
rect 402 792 406 796
rect 732 800 736 804
rect 874 800 878 804
rect 1014 800 1018 804
rect 1159 800 1163 804
rect 1304 800 1308 804
rect 1449 800 1453 804
rect 402 784 406 788
rect 518 786 522 790
rect 148 756 152 760
rect 148 748 152 752
rect 732 749 736 753
rect 874 749 878 753
rect 1014 749 1018 753
rect 1159 749 1163 753
rect 1304 749 1308 753
rect 1449 749 1453 753
rect -1144 727 -1140 731
rect -1144 719 -1140 723
rect -817 727 -813 731
rect -1250 709 -1246 713
rect -817 719 -813 723
rect -485 726 -481 730
rect -1250 701 -1246 705
rect -923 709 -919 713
rect -485 718 -481 722
rect -158 726 -154 730
rect -923 701 -919 705
rect -591 708 -587 712
rect -158 718 -154 722
rect 57 722 61 726
rect -591 700 -587 704
rect -264 708 -260 712
rect 57 714 61 718
rect 244 722 248 726
rect 244 714 248 718
rect 361 715 365 719
rect -264 700 -260 704
rect 148 700 152 704
rect 361 707 365 711
rect 148 692 152 696
rect 361 699 365 703
rect 439 707 443 711
rect 457 700 461 704
rect -1329 654 -1325 658
rect -1278 654 -1274 658
rect -1250 662 -1246 666
rect -1250 654 -1246 658
rect -1144 662 -1140 666
rect -1144 654 -1140 658
rect -1001 654 -997 658
rect -951 654 -947 658
rect -923 662 -919 666
rect -923 654 -919 658
rect -817 662 -813 666
rect -817 654 -813 658
rect -670 653 -666 657
rect -619 653 -615 657
rect -591 661 -587 665
rect -591 653 -587 657
rect -485 661 -481 665
rect -485 653 -481 657
rect -342 653 -338 657
rect -292 653 -288 657
rect -264 661 -260 665
rect -264 653 -260 657
rect -158 661 -154 665
rect -158 653 -154 657
rect 639 669 643 673
rect 639 661 643 665
rect 45 642 49 646
rect 45 634 49 638
rect 132 638 136 642
rect 280 629 284 633
rect 548 635 552 639
rect 280 621 284 625
rect 548 627 552 631
rect 735 635 739 639
rect 735 627 739 631
rect 639 613 643 617
rect 639 605 643 609
rect 189 595 193 599
rect 189 587 193 591
rect 376 595 380 599
rect 376 587 380 591
rect 280 573 284 577
rect 280 565 284 569
rect 535 531 539 535
rect 535 523 539 527
rect 622 527 626 531
rect -1144 513 -1140 517
rect -1144 505 -1140 509
rect -817 513 -813 517
rect -1250 495 -1246 499
rect -817 505 -813 509
rect -485 512 -481 516
rect -1250 487 -1246 491
rect -923 495 -919 499
rect -485 504 -481 508
rect -158 512 -154 516
rect -923 487 -919 491
rect -591 494 -587 498
rect -158 504 -154 508
rect -591 486 -587 490
rect -264 494 -260 498
rect 148 502 152 506
rect -264 486 -260 490
rect 148 494 152 498
rect 366 480 370 484
rect -1329 440 -1325 444
rect -1278 440 -1274 444
rect -1250 448 -1246 452
rect -1250 440 -1246 444
rect -1144 448 -1140 452
rect -1144 440 -1140 444
rect -1001 440 -997 444
rect -951 440 -947 444
rect -923 448 -919 452
rect -923 440 -919 444
rect -817 448 -813 452
rect -817 440 -813 444
rect -670 439 -666 443
rect -619 439 -615 443
rect -591 447 -587 451
rect -591 439 -587 443
rect -485 447 -481 451
rect 57 468 61 472
rect 57 460 61 464
rect 244 468 248 472
rect 366 472 370 476
rect 535 478 539 482
rect 244 460 248 464
rect 366 464 370 468
rect 366 456 370 460
rect 454 464 458 468
rect 472 462 476 466
rect 535 470 539 474
rect 682 494 686 498
rect 682 486 686 490
rect 682 478 686 482
rect 535 462 539 466
rect 631 463 635 467
rect -485 439 -481 443
rect -342 439 -338 443
rect -292 439 -288 443
rect -264 447 -260 451
rect -264 439 -260 443
rect -158 447 -154 451
rect -158 439 -154 443
rect 148 446 152 450
rect 682 470 686 474
rect 819 474 823 478
rect 148 438 152 442
rect 712 410 716 414
rect 781 411 785 415
rect 712 402 716 406
rect 799 406 803 410
rect 45 388 49 392
rect 45 380 49 384
rect 132 384 136 388
rect 294 367 298 371
rect 294 359 298 363
rect 430 369 434 373
rect 294 351 298 355
rect 294 343 298 347
rect 367 351 371 355
rect 386 350 390 354
rect 430 361 434 365
rect 576 366 580 370
rect 430 353 434 357
rect 294 335 298 339
rect 375 337 379 341
rect 430 345 434 349
rect 518 353 522 357
rect 536 351 540 355
rect 576 358 580 362
rect 576 350 580 354
rect 654 350 658 354
rect 672 351 676 355
rect 722 346 726 350
rect 722 338 726 342
rect 722 330 726 334
rect 149 320 153 324
rect 722 322 726 326
rect 877 330 881 334
rect 149 312 153 316
rect 722 314 726 318
rect 58 286 62 290
rect -1144 274 -1140 278
rect -1144 266 -1140 270
rect -817 274 -813 278
rect -1250 256 -1246 260
rect -817 266 -813 270
rect -485 273 -481 277
rect -1250 248 -1246 252
rect -923 256 -919 260
rect -485 265 -481 269
rect -158 273 -154 277
rect 58 278 62 282
rect 245 286 249 290
rect 245 278 249 282
rect -923 248 -919 252
rect -591 255 -587 259
rect -158 265 -154 269
rect -591 247 -587 251
rect -264 255 -260 259
rect 149 264 153 268
rect 149 256 153 260
rect -264 247 -260 251
rect 472 251 476 255
rect 472 243 476 247
rect 1097 248 1101 252
rect 1097 240 1101 244
rect -1329 201 -1325 205
rect -1278 201 -1274 205
rect -1250 209 -1246 213
rect -1250 201 -1246 205
rect -1144 209 -1140 213
rect -1144 201 -1140 205
rect -1001 201 -997 205
rect -951 201 -947 205
rect -923 209 -919 213
rect -923 201 -919 205
rect -817 209 -813 213
rect -817 201 -813 205
rect -670 200 -666 204
rect -619 200 -615 204
rect -591 208 -587 212
rect -591 200 -587 204
rect -485 208 -481 212
rect -485 200 -481 204
rect -342 200 -338 204
rect -292 200 -288 204
rect -264 208 -260 212
rect -264 200 -260 204
rect -158 208 -154 212
rect 381 217 385 221
rect -158 200 -154 204
rect 46 206 50 210
rect 46 198 50 202
rect 133 202 137 206
rect 381 209 385 213
rect 568 217 572 221
rect 568 209 572 213
rect 472 195 476 199
rect 693 198 697 202
rect 472 187 476 191
rect 693 190 697 194
rect 839 210 843 214
rect 839 202 843 206
rect 926 206 930 210
rect 1006 214 1010 218
rect 1006 206 1010 210
rect 1193 214 1197 218
rect 693 182 697 186
rect 789 183 793 187
rect 1193 206 1197 210
rect 1097 192 1101 196
rect 1097 184 1101 188
rect 150 137 154 141
rect 150 129 154 133
rect 375 127 379 131
rect 375 119 379 123
rect 375 111 379 115
rect 512 129 516 133
rect 512 121 516 125
rect 59 103 63 107
rect 59 95 63 99
rect 246 103 250 107
rect -1144 87 -1140 91
rect -1144 79 -1140 83
rect -817 87 -813 91
rect -1250 69 -1246 73
rect -817 79 -813 83
rect -485 86 -481 90
rect -1250 61 -1246 65
rect -923 69 -919 73
rect -485 78 -481 82
rect -158 86 -154 90
rect 246 95 250 99
rect 375 103 379 107
rect 446 111 450 115
rect 375 95 379 99
rect 446 102 450 106
rect 471 103 475 107
rect 512 113 516 117
rect 512 105 516 109
rect 585 113 589 117
rect 604 112 608 116
rect 640 121 644 125
rect 640 113 644 117
rect 849 125 853 129
rect 849 117 853 121
rect -923 61 -919 65
rect -591 68 -587 72
rect -158 78 -154 82
rect 150 81 154 85
rect 375 87 379 91
rect 446 94 450 98
rect 512 97 516 101
rect 594 102 598 106
rect 640 105 644 109
rect 640 97 644 101
rect 728 105 732 109
rect 746 103 750 107
rect 849 109 853 113
rect 849 101 853 105
rect 849 93 853 97
rect 1035 101 1039 105
rect 849 85 853 89
rect -591 60 -587 64
rect -264 68 -260 72
rect 150 73 154 77
rect -264 60 -260 64
rect -1329 14 -1325 18
rect -1278 14 -1274 18
rect -1250 22 -1246 26
rect -1250 14 -1246 18
rect -1144 22 -1140 26
rect -1144 14 -1140 18
rect -1001 14 -997 18
rect -951 14 -947 18
rect -923 22 -919 26
rect -923 14 -919 18
rect -817 22 -813 26
rect -817 14 -813 18
rect -670 13 -666 17
rect -619 13 -615 17
rect -591 21 -587 25
rect -591 13 -587 17
rect -485 21 -481 25
rect -485 13 -481 17
rect -342 13 -338 17
rect -292 13 -288 17
rect -264 21 -260 25
rect -264 13 -260 17
rect -158 21 -154 25
rect 47 23 51 27
rect -158 13 -154 17
rect 47 15 51 19
rect 134 19 138 23
<< ndcontact >>
rect 655 1313 659 1333
rect 663 1313 667 1333
rect 671 1313 675 1333
rect 720 1313 724 1333
rect 728 1313 732 1333
rect 736 1313 740 1333
rect 797 1313 801 1333
rect 805 1313 809 1333
rect 813 1313 817 1333
rect 862 1313 866 1333
rect 870 1313 874 1333
rect 878 1313 882 1333
rect 937 1313 941 1333
rect 945 1313 949 1333
rect 953 1313 957 1333
rect 1002 1313 1006 1333
rect 1010 1313 1014 1333
rect 1018 1313 1022 1333
rect 1082 1313 1086 1333
rect 1090 1313 1094 1333
rect 1098 1313 1102 1333
rect 1147 1313 1151 1333
rect 1155 1313 1159 1333
rect 1163 1313 1167 1333
rect 1227 1313 1231 1333
rect 1235 1313 1239 1333
rect 1243 1313 1247 1333
rect 1292 1313 1296 1333
rect 1300 1313 1304 1333
rect 1308 1313 1312 1333
rect 1372 1313 1376 1333
rect 1380 1313 1384 1333
rect 1388 1313 1392 1333
rect 1437 1313 1441 1333
rect 1445 1313 1449 1333
rect 1453 1313 1457 1333
rect 673 1207 677 1227
rect 681 1207 685 1227
rect 689 1207 693 1227
rect 720 1207 724 1227
rect 728 1207 732 1227
rect 736 1207 740 1227
rect 815 1207 819 1227
rect 823 1207 827 1227
rect 831 1207 835 1227
rect 862 1207 866 1227
rect 870 1207 874 1227
rect 878 1207 882 1227
rect 955 1207 959 1227
rect 963 1207 967 1227
rect 971 1207 975 1227
rect 1002 1207 1006 1227
rect 1010 1207 1014 1227
rect 1018 1207 1022 1227
rect 1100 1207 1104 1227
rect 1108 1207 1112 1227
rect 1116 1207 1120 1227
rect 1147 1207 1151 1227
rect 1155 1207 1159 1227
rect 1163 1207 1167 1227
rect 1245 1207 1249 1227
rect 1253 1207 1257 1227
rect 1261 1207 1265 1227
rect 1292 1207 1296 1227
rect 1300 1207 1304 1227
rect 1308 1207 1312 1227
rect 1390 1207 1394 1227
rect 1398 1207 1402 1227
rect 1406 1207 1410 1227
rect 1437 1207 1441 1227
rect 1445 1207 1449 1227
rect 1453 1207 1457 1227
rect -432 1130 -412 1134
rect -105 1130 -85 1134
rect 739 1134 749 1138
rect 881 1134 891 1138
rect 1021 1134 1031 1138
rect 1166 1134 1176 1138
rect 1311 1134 1321 1138
rect 1456 1134 1466 1138
rect -432 1122 -412 1126
rect -538 1112 -518 1116
rect 739 1126 749 1130
rect 881 1126 891 1130
rect 1021 1126 1031 1130
rect 1166 1126 1176 1130
rect 1311 1126 1321 1130
rect 1456 1126 1466 1130
rect -105 1122 -85 1126
rect -432 1114 -412 1118
rect -211 1112 -191 1116
rect -105 1114 -85 1118
rect -538 1104 -518 1108
rect -211 1104 -191 1108
rect -538 1096 -518 1100
rect -211 1096 -191 1100
rect -538 1065 -518 1069
rect -432 1065 -412 1069
rect 739 1084 749 1088
rect 881 1084 891 1088
rect 1021 1084 1031 1088
rect 1166 1084 1176 1088
rect 1311 1084 1321 1088
rect 1456 1084 1466 1088
rect 739 1076 749 1080
rect 881 1076 891 1080
rect 1021 1076 1031 1080
rect 1166 1076 1176 1080
rect 1311 1076 1321 1080
rect 1456 1076 1466 1080
rect -538 1057 -518 1061
rect -670 1040 -666 1050
rect -662 1040 -658 1050
rect -619 1040 -615 1050
rect -611 1040 -607 1050
rect -432 1057 -412 1061
rect -538 1049 -518 1053
rect -432 1049 -412 1053
rect -211 1065 -191 1069
rect -105 1065 -85 1069
rect -211 1057 -191 1061
rect -342 1040 -338 1050
rect -334 1040 -330 1050
rect -292 1040 -288 1050
rect -284 1040 -280 1050
rect -105 1057 -85 1061
rect -211 1049 -191 1053
rect -105 1049 -85 1053
rect 452 1028 472 1032
rect 452 1020 472 1024
rect 452 1012 472 1016
rect 361 994 381 998
rect 548 994 568 998
rect 361 986 381 990
rect 548 986 568 990
rect 655 986 659 1006
rect 663 986 667 1006
rect 671 986 675 1006
rect 720 986 724 1006
rect 728 986 732 1006
rect 736 986 740 1006
rect 797 986 801 1006
rect 805 986 809 1006
rect 813 986 817 1006
rect 862 986 866 1006
rect 870 986 874 1006
rect 878 986 882 1006
rect 937 986 941 1006
rect 945 986 949 1006
rect 953 986 957 1006
rect 1002 986 1006 1006
rect 1010 986 1014 1006
rect 1018 986 1022 1006
rect 1082 986 1086 1006
rect 1090 986 1094 1006
rect 1098 986 1102 1006
rect 1147 986 1151 1006
rect 1155 986 1159 1006
rect 1163 986 1167 1006
rect 1227 986 1231 1006
rect 1235 986 1239 1006
rect 1243 986 1247 1006
rect 1292 986 1296 1006
rect 1300 986 1304 1006
rect 1308 986 1312 1006
rect 1372 986 1376 1006
rect 1380 986 1384 1006
rect 1388 986 1392 1006
rect 1437 986 1441 1006
rect 1445 986 1449 1006
rect 1453 986 1457 1006
rect 361 978 381 982
rect 548 978 568 982
rect -1092 970 -1072 974
rect -765 970 -745 974
rect -1092 962 -1072 966
rect -1198 952 -1178 956
rect -765 962 -745 966
rect -433 966 -413 970
rect -1092 954 -1072 958
rect -871 952 -851 956
rect -765 954 -745 958
rect -106 966 -86 970
rect 452 972 472 976
rect -433 958 -413 962
rect -1198 944 -1178 948
rect -871 944 -851 948
rect -539 948 -519 952
rect -106 958 -86 962
rect 452 964 472 968
rect 452 956 472 960
rect -433 950 -413 954
rect -1198 936 -1178 940
rect -871 936 -851 940
rect -212 948 -192 952
rect -106 950 -86 954
rect -539 940 -519 944
rect -212 940 -192 944
rect -539 932 -519 936
rect 201 940 221 944
rect -212 932 -192 936
rect 201 932 221 936
rect 201 924 221 928
rect -1198 905 -1178 909
rect -1092 905 -1072 909
rect -1198 897 -1178 901
rect -1330 880 -1326 890
rect -1322 880 -1318 890
rect -1279 880 -1275 890
rect -1271 880 -1267 890
rect -1092 897 -1072 901
rect -1198 889 -1178 893
rect -1092 889 -1072 893
rect -871 905 -851 909
rect -765 905 -745 909
rect -871 897 -851 901
rect -1002 880 -998 890
rect -994 880 -990 890
rect -952 880 -948 890
rect -944 880 -940 890
rect -765 897 -745 901
rect -871 889 -851 893
rect -765 889 -745 893
rect -539 901 -519 905
rect -433 901 -413 905
rect -539 893 -519 897
rect -671 876 -667 886
rect -663 876 -659 886
rect -620 876 -616 886
rect -612 876 -608 886
rect -433 893 -413 897
rect -539 885 -519 889
rect -433 885 -413 889
rect -212 901 -192 905
rect -106 901 -86 905
rect 110 906 130 910
rect -212 893 -192 897
rect -343 876 -339 886
rect -335 876 -331 886
rect -293 876 -289 886
rect -285 876 -281 886
rect -106 893 -86 897
rect 297 906 317 910
rect 110 898 130 902
rect 297 898 317 902
rect 110 890 130 894
rect 297 890 317 894
rect -212 885 -192 889
rect -106 885 -86 889
rect 201 884 221 888
rect 401 887 421 891
rect 201 876 221 880
rect 401 879 421 883
rect 538 886 548 890
rect 201 868 221 872
rect 401 871 421 875
rect 441 866 445 876
rect 449 866 453 876
rect 538 878 548 882
rect 673 880 677 900
rect 681 880 685 900
rect 689 880 693 900
rect 720 880 724 900
rect 728 880 732 900
rect 736 880 740 900
rect 815 880 819 900
rect 823 880 827 900
rect 831 880 835 900
rect 862 880 866 900
rect 870 880 874 900
rect 878 880 882 900
rect 955 880 959 900
rect 963 880 967 900
rect 971 880 975 900
rect 1002 880 1006 900
rect 1010 880 1014 900
rect 1018 880 1022 900
rect 1100 880 1104 900
rect 1108 880 1112 900
rect 1116 880 1120 900
rect 1147 880 1151 900
rect 1155 880 1159 900
rect 1163 880 1167 900
rect 1245 880 1249 900
rect 1253 880 1257 900
rect 1261 880 1265 900
rect 1292 880 1296 900
rect 1300 880 1304 900
rect 1308 880 1312 900
rect 1390 880 1394 900
rect 1398 880 1402 900
rect 1406 880 1410 900
rect 1437 880 1441 900
rect 1445 880 1449 900
rect 1453 880 1457 900
rect 538 870 548 874
rect 569 866 573 876
rect 577 866 581 876
rect 92 826 112 830
rect 92 818 112 822
rect 92 810 112 814
rect 132 805 136 815
rect 140 805 144 815
rect 324 801 344 805
rect 324 793 344 797
rect 487 804 497 808
rect 487 796 497 800
rect 739 807 749 811
rect 881 807 891 811
rect 1021 807 1031 811
rect 1166 807 1176 811
rect 1311 807 1321 811
rect 1456 807 1466 811
rect 739 799 749 803
rect 881 799 891 803
rect 1021 799 1031 803
rect 1166 799 1176 803
rect 1311 799 1321 803
rect 1456 799 1466 803
rect 324 785 344 789
rect 364 780 368 790
rect 372 780 376 790
rect 487 788 497 792
rect 487 780 497 784
rect 517 773 521 783
rect 525 773 529 783
rect 200 760 220 764
rect 200 752 220 756
rect 739 756 749 760
rect 881 756 891 760
rect 1021 756 1031 760
rect 1166 756 1176 760
rect 1311 756 1321 760
rect 1456 756 1466 760
rect 739 748 749 752
rect 881 748 891 752
rect 1021 748 1031 752
rect 1166 748 1176 752
rect 1311 748 1321 752
rect 1456 748 1466 752
rect 200 744 220 748
rect -1092 731 -1072 735
rect -765 731 -745 735
rect -1092 723 -1072 727
rect -1198 713 -1178 717
rect -765 723 -745 727
rect -433 730 -413 734
rect -1092 715 -1072 719
rect -871 713 -851 717
rect -765 715 -745 719
rect -106 730 -86 734
rect -433 722 -413 726
rect -1198 705 -1178 709
rect -871 705 -851 709
rect -539 712 -519 716
rect -106 722 -86 726
rect 109 726 129 730
rect -433 714 -413 718
rect -1198 697 -1178 701
rect -871 697 -851 701
rect -212 712 -192 716
rect -106 714 -86 718
rect 296 726 316 730
rect 109 718 129 722
rect 296 718 316 722
rect 406 719 436 723
rect 109 710 129 714
rect 296 710 316 714
rect -539 704 -519 708
rect -212 704 -192 708
rect -539 696 -519 700
rect 200 704 220 708
rect 406 711 436 715
rect -212 696 -192 700
rect 200 696 220 700
rect 406 703 436 707
rect 406 695 436 699
rect 200 688 220 692
rect 456 687 460 697
rect 464 687 468 697
rect -1198 666 -1178 670
rect -1092 666 -1072 670
rect -1198 658 -1178 662
rect -1330 641 -1326 651
rect -1322 641 -1318 651
rect -1279 641 -1275 651
rect -1271 641 -1267 651
rect -1092 658 -1072 662
rect -1198 650 -1178 654
rect -1092 650 -1072 654
rect -871 666 -851 670
rect -765 666 -745 670
rect -871 658 -851 662
rect -1002 641 -998 651
rect -994 641 -990 651
rect -952 641 -948 651
rect -944 641 -940 651
rect -765 658 -745 662
rect -871 650 -851 654
rect -765 650 -745 654
rect -539 665 -519 669
rect -433 665 -413 669
rect -539 657 -519 661
rect -671 640 -667 650
rect -663 640 -659 650
rect -620 640 -616 650
rect -612 640 -608 650
rect -433 657 -413 661
rect -539 649 -519 653
rect -433 649 -413 653
rect -212 665 -192 669
rect -106 665 -86 669
rect -212 657 -192 661
rect -343 640 -339 650
rect -335 640 -331 650
rect -293 640 -289 650
rect -285 640 -281 650
rect -106 657 -86 661
rect -212 649 -192 653
rect -106 649 -86 653
rect 691 673 711 677
rect 691 665 711 669
rect 691 657 711 661
rect 91 646 111 650
rect 91 638 111 642
rect 91 630 111 634
rect 131 625 135 635
rect 139 625 143 635
rect 332 633 352 637
rect 600 639 620 643
rect 332 625 352 629
rect 787 639 807 643
rect 600 631 620 635
rect 787 631 807 635
rect 600 623 620 627
rect 787 623 807 627
rect 332 617 352 621
rect 691 617 711 621
rect 691 609 711 613
rect 241 599 261 603
rect 428 599 448 603
rect 691 601 711 605
rect 241 591 261 595
rect 428 591 448 595
rect 241 583 261 587
rect 428 583 448 587
rect 332 577 352 581
rect 332 569 352 573
rect 332 561 352 565
rect 581 535 601 539
rect 581 527 601 531
rect -1092 517 -1072 521
rect -765 517 -745 521
rect -1092 509 -1072 513
rect -1198 499 -1178 503
rect -765 509 -745 513
rect -433 516 -413 520
rect -1092 501 -1072 505
rect -871 499 -851 503
rect -765 501 -745 505
rect -106 516 -86 520
rect 581 519 601 523
rect 621 514 625 524
rect 629 514 633 524
rect -433 508 -413 512
rect -1198 491 -1178 495
rect -871 491 -851 495
rect -539 498 -519 502
rect -106 508 -86 512
rect -433 500 -413 504
rect -1198 483 -1178 487
rect -871 483 -851 487
rect -212 498 -192 502
rect -106 500 -86 504
rect 200 506 220 510
rect -539 490 -519 494
rect 200 498 220 502
rect -212 490 -192 494
rect 200 490 220 494
rect -539 482 -519 486
rect -212 482 -192 486
rect 411 484 451 488
rect -1198 452 -1178 456
rect -1092 452 -1072 456
rect -1198 444 -1178 448
rect -1330 427 -1326 437
rect -1322 427 -1318 437
rect -1279 427 -1275 437
rect -1271 427 -1267 437
rect -1092 444 -1072 448
rect -1198 436 -1178 440
rect -1092 436 -1072 440
rect -871 452 -851 456
rect -765 452 -745 456
rect -871 444 -851 448
rect -1002 427 -998 437
rect -994 427 -990 437
rect -952 427 -948 437
rect -944 427 -940 437
rect -765 444 -745 448
rect -871 436 -851 440
rect -765 436 -745 440
rect -539 451 -519 455
rect -433 451 -413 455
rect 109 472 129 476
rect 296 472 316 476
rect 411 476 451 480
rect 580 482 610 486
rect 109 464 129 468
rect 296 464 316 468
rect 411 468 451 472
rect 109 456 129 460
rect 296 456 316 460
rect 411 460 451 464
rect 580 474 610 478
rect 787 498 797 502
rect 787 490 797 494
rect 787 482 797 486
rect 580 466 610 470
rect -539 443 -519 447
rect -671 426 -667 436
rect -663 426 -659 436
rect -620 426 -616 436
rect -612 426 -608 436
rect -433 443 -413 447
rect -539 435 -519 439
rect -433 435 -413 439
rect -212 451 -192 455
rect -106 451 -86 455
rect -212 443 -192 447
rect -343 426 -339 436
rect -335 426 -331 436
rect -293 426 -289 436
rect -285 426 -281 436
rect -106 443 -86 447
rect 200 450 220 454
rect 411 452 451 456
rect 471 449 475 459
rect 479 449 483 459
rect 580 458 610 462
rect 787 474 797 478
rect 787 466 797 470
rect 818 461 822 471
rect 826 461 830 471
rect 630 450 634 460
rect 638 450 642 460
rect -212 435 -192 439
rect -106 435 -86 439
rect 200 442 220 446
rect 200 434 220 438
rect 758 414 778 418
rect 758 406 778 410
rect 758 398 778 402
rect 91 392 111 396
rect 91 384 111 388
rect 798 393 802 403
rect 806 393 810 403
rect 91 376 111 380
rect 131 371 135 381
rect 139 371 143 381
rect 339 371 364 375
rect 339 363 364 367
rect 475 373 515 377
rect 339 355 364 359
rect 339 347 364 351
rect 475 365 515 369
rect 621 370 651 374
rect 475 357 515 361
rect 339 339 364 343
rect 385 337 389 347
rect 393 337 397 347
rect 475 349 515 353
rect 621 362 651 366
rect 621 354 651 358
rect 475 341 515 345
rect 535 338 539 348
rect 543 338 547 348
rect 621 346 651 350
rect 671 338 675 348
rect 679 338 683 348
rect 847 350 857 354
rect 847 342 857 346
rect 339 331 364 335
rect 847 334 857 338
rect 201 324 221 328
rect 847 326 857 330
rect 201 316 221 320
rect 847 318 857 322
rect 876 317 880 327
rect 884 317 888 327
rect 201 308 221 312
rect 847 310 857 314
rect 110 290 130 294
rect -1092 278 -1072 282
rect -765 278 -745 282
rect -1092 270 -1072 274
rect -1198 260 -1178 264
rect -765 270 -745 274
rect -433 277 -413 281
rect -1092 262 -1072 266
rect -871 260 -851 264
rect -765 262 -745 266
rect -106 277 -86 281
rect 297 290 317 294
rect 110 282 130 286
rect 297 282 317 286
rect 110 274 130 278
rect 297 274 317 278
rect -433 269 -413 273
rect -1198 252 -1178 256
rect -871 252 -851 256
rect -539 259 -519 263
rect -106 269 -86 273
rect -433 261 -413 265
rect -1198 244 -1178 248
rect -871 244 -851 248
rect -212 259 -192 263
rect -106 261 -86 265
rect 201 268 221 272
rect 201 260 221 264
rect -539 251 -519 255
rect -212 251 -192 255
rect 201 252 221 256
rect 524 255 544 259
rect -539 243 -519 247
rect -212 243 -192 247
rect 524 247 544 251
rect 1149 252 1169 256
rect 524 239 544 243
rect 1149 244 1169 248
rect -1198 213 -1178 217
rect -1092 213 -1072 217
rect -1198 205 -1178 209
rect -1330 188 -1326 198
rect -1322 188 -1318 198
rect -1279 188 -1275 198
rect -1271 188 -1267 198
rect -1092 205 -1072 209
rect -1198 197 -1178 201
rect -1092 197 -1072 201
rect -871 213 -851 217
rect -765 213 -745 217
rect -871 205 -851 209
rect -1002 188 -998 198
rect -994 188 -990 198
rect -952 188 -948 198
rect -944 188 -940 198
rect -765 205 -745 209
rect -871 197 -851 201
rect -765 197 -745 201
rect -539 212 -519 216
rect -433 212 -413 216
rect -539 204 -519 208
rect -671 187 -667 197
rect -663 187 -659 197
rect -620 187 -616 197
rect -612 187 -608 197
rect -433 204 -413 208
rect -539 196 -519 200
rect -433 196 -413 200
rect -212 212 -192 216
rect -106 212 -86 216
rect 433 221 453 225
rect -212 204 -192 208
rect -343 187 -339 197
rect -335 187 -331 197
rect -293 187 -289 197
rect -285 187 -281 197
rect -106 204 -86 208
rect 92 210 112 214
rect -212 196 -192 200
rect -106 196 -86 200
rect 92 202 112 206
rect 620 221 640 225
rect 1149 236 1169 240
rect 433 213 453 217
rect 620 213 640 217
rect 433 205 453 209
rect 620 205 640 209
rect 92 194 112 198
rect 132 189 136 199
rect 140 189 144 199
rect 524 199 544 203
rect 738 202 768 206
rect 524 191 544 195
rect 738 194 768 198
rect 885 214 905 218
rect 885 206 905 210
rect 1058 218 1078 222
rect 1245 218 1265 222
rect 1058 210 1078 214
rect 885 198 905 202
rect 524 183 544 187
rect 738 186 768 190
rect 738 178 768 182
rect 925 193 929 203
rect 933 193 937 203
rect 1245 210 1265 214
rect 1058 202 1078 206
rect 1245 202 1265 206
rect 1149 196 1169 200
rect 1149 188 1169 192
rect 1149 180 1169 184
rect 788 170 792 180
rect 796 170 800 180
rect 202 141 222 145
rect 202 133 222 137
rect 202 125 222 129
rect 413 131 443 135
rect 413 123 443 127
rect 413 115 443 119
rect 557 133 582 137
rect 557 125 582 129
rect 111 107 131 111
rect 298 107 318 111
rect 111 99 131 103
rect -1092 91 -1072 95
rect -765 91 -745 95
rect -1092 83 -1072 87
rect -1198 73 -1178 77
rect -765 83 -745 87
rect -433 90 -413 94
rect -1092 75 -1072 79
rect -871 73 -851 77
rect -765 75 -745 79
rect -106 90 -86 94
rect 413 107 443 111
rect 298 99 318 103
rect 111 91 131 95
rect 413 99 443 103
rect 557 117 582 121
rect 557 109 582 113
rect 685 125 725 129
rect 685 117 725 121
rect 996 129 1006 133
rect 996 121 1006 125
rect 298 91 318 95
rect -433 82 -413 86
rect -1198 65 -1178 69
rect -871 65 -851 69
rect -539 72 -519 76
rect -106 82 -86 86
rect 202 85 222 89
rect 413 91 443 95
rect 470 90 474 100
rect 478 90 482 100
rect 557 101 582 105
rect 603 99 607 109
rect 611 99 615 109
rect 685 109 725 113
rect 557 93 582 97
rect 685 101 725 105
rect 996 113 1006 117
rect 996 105 1006 109
rect 685 93 725 97
rect 745 90 749 100
rect 753 90 757 100
rect 996 97 1006 101
rect 413 83 443 87
rect 996 89 1006 93
rect 1034 88 1038 98
rect 1042 88 1046 98
rect -433 74 -413 78
rect -1198 57 -1178 61
rect -871 57 -851 61
rect -212 72 -192 76
rect -106 74 -86 78
rect 996 81 1006 85
rect 202 77 222 81
rect 202 69 222 73
rect -539 64 -519 68
rect -212 64 -192 68
rect -539 56 -519 60
rect -212 56 -192 60
rect -1198 26 -1178 30
rect -1092 26 -1072 30
rect -1198 18 -1178 22
rect -1330 1 -1326 11
rect -1322 1 -1318 11
rect -1279 1 -1275 11
rect -1271 1 -1267 11
rect -1092 18 -1072 22
rect -1198 10 -1178 14
rect -1092 10 -1072 14
rect -871 26 -851 30
rect -765 26 -745 30
rect -871 18 -851 22
rect -1002 1 -998 11
rect -994 1 -990 11
rect -952 1 -948 11
rect -944 1 -940 11
rect -765 18 -745 22
rect -871 10 -851 14
rect -765 10 -745 14
rect -539 25 -519 29
rect -433 25 -413 29
rect -539 17 -519 21
rect -671 0 -667 10
rect -663 0 -659 10
rect -620 0 -616 10
rect -612 0 -608 10
rect -433 17 -413 21
rect -539 9 -519 13
rect -433 9 -413 13
rect -212 25 -192 29
rect -106 25 -86 29
rect 93 27 113 31
rect -212 17 -192 21
rect -343 0 -339 10
rect -335 0 -331 10
rect -293 0 -289 10
rect -285 0 -281 10
rect -106 17 -86 21
rect 93 19 113 23
rect -212 9 -192 13
rect -106 9 -86 13
rect 93 11 113 15
rect 133 6 137 16
rect 141 6 145 16
<< pdcontact >>
rect 655 1277 659 1297
rect 663 1277 667 1297
rect 671 1277 675 1297
rect 720 1277 724 1297
rect 728 1277 732 1297
rect 736 1277 740 1297
rect 797 1277 801 1297
rect 805 1277 809 1297
rect 813 1277 817 1297
rect 862 1277 866 1297
rect 870 1277 874 1297
rect 878 1277 882 1297
rect 937 1277 941 1297
rect 945 1277 949 1297
rect 953 1277 957 1297
rect 1002 1277 1006 1297
rect 1010 1277 1014 1297
rect 1018 1277 1022 1297
rect 1082 1277 1086 1297
rect 1090 1277 1094 1297
rect 1098 1277 1102 1297
rect 1147 1277 1151 1297
rect 1155 1277 1159 1297
rect 1163 1277 1167 1297
rect 1227 1277 1231 1297
rect 1235 1277 1239 1297
rect 1243 1277 1247 1297
rect 1292 1277 1296 1297
rect 1300 1277 1304 1297
rect 1308 1277 1312 1297
rect 1372 1277 1376 1297
rect 1380 1277 1384 1297
rect 1388 1277 1392 1297
rect 1437 1277 1441 1297
rect 1445 1277 1449 1297
rect 1453 1277 1457 1297
rect 673 1171 677 1191
rect 681 1171 685 1191
rect 689 1171 693 1191
rect 720 1171 724 1191
rect 728 1171 732 1191
rect 736 1171 740 1191
rect 815 1171 819 1191
rect 823 1171 827 1191
rect 831 1171 835 1191
rect 862 1171 866 1191
rect 870 1171 874 1191
rect 878 1171 882 1191
rect 955 1171 959 1191
rect 963 1171 967 1191
rect 971 1171 975 1191
rect 1002 1171 1006 1191
rect 1010 1171 1014 1191
rect 1018 1171 1022 1191
rect 1100 1171 1104 1191
rect 1108 1171 1112 1191
rect 1116 1171 1120 1191
rect 1147 1171 1151 1191
rect 1155 1171 1159 1191
rect 1163 1171 1167 1191
rect 1245 1171 1249 1191
rect 1253 1171 1257 1191
rect 1261 1171 1265 1191
rect 1292 1171 1296 1191
rect 1300 1171 1304 1191
rect 1308 1171 1312 1191
rect 1390 1171 1394 1191
rect 1398 1171 1402 1191
rect 1406 1171 1410 1191
rect 1437 1171 1441 1191
rect 1445 1171 1449 1191
rect 1453 1171 1457 1191
rect 705 1134 725 1138
rect -468 1130 -448 1134
rect -141 1130 -121 1134
rect -468 1122 -448 1126
rect 847 1134 867 1138
rect 987 1134 1007 1138
rect 1132 1134 1152 1138
rect 1277 1134 1297 1138
rect 1422 1134 1442 1138
rect -141 1122 -121 1126
rect -574 1112 -554 1116
rect -468 1114 -448 1118
rect 705 1126 725 1130
rect 847 1126 867 1130
rect 987 1126 1007 1130
rect 1132 1126 1152 1130
rect 1277 1126 1297 1130
rect 1422 1126 1442 1130
rect -247 1112 -227 1116
rect -574 1104 -554 1108
rect -141 1114 -121 1118
rect -247 1104 -227 1108
rect -574 1096 -554 1100
rect -247 1096 -227 1100
rect 705 1084 725 1088
rect -670 1064 -666 1084
rect -662 1064 -658 1084
rect -619 1064 -615 1084
rect -611 1064 -607 1084
rect -574 1065 -554 1069
rect -468 1065 -448 1069
rect -574 1057 -554 1061
rect -342 1064 -338 1084
rect -334 1064 -330 1084
rect -292 1064 -288 1084
rect -284 1064 -280 1084
rect 847 1084 867 1088
rect 987 1084 1007 1088
rect 1132 1084 1152 1088
rect 1277 1084 1297 1088
rect 1422 1084 1442 1088
rect 705 1076 725 1080
rect 847 1076 867 1080
rect 987 1076 1007 1080
rect 1132 1076 1152 1080
rect 1277 1076 1297 1080
rect 1422 1076 1442 1080
rect -247 1065 -227 1069
rect -468 1057 -448 1061
rect -574 1049 -554 1053
rect -468 1049 -448 1053
rect -141 1065 -121 1069
rect -247 1057 -227 1061
rect -141 1057 -121 1061
rect -247 1049 -227 1053
rect -141 1049 -121 1053
rect 416 1028 436 1032
rect 416 1020 436 1024
rect 416 1012 436 1016
rect 325 994 345 998
rect 512 994 532 998
rect 325 986 345 990
rect 512 986 532 990
rect 325 978 345 982
rect 512 978 532 982
rect -1128 970 -1108 974
rect -801 970 -781 974
rect -1128 962 -1108 966
rect 416 972 436 976
rect -801 962 -781 966
rect -1234 952 -1214 956
rect -1128 954 -1108 958
rect -469 966 -449 970
rect -142 966 -122 970
rect -907 952 -887 956
rect -1234 944 -1214 948
rect -801 954 -781 958
rect -469 958 -449 962
rect 416 964 436 968
rect -142 958 -122 962
rect -907 944 -887 948
rect -1234 936 -1214 940
rect -575 948 -555 952
rect -469 950 -449 954
rect 416 956 436 960
rect -248 948 -228 952
rect -907 936 -887 940
rect -575 940 -555 944
rect -142 950 -122 954
rect 655 950 659 970
rect 663 950 667 970
rect 671 950 675 970
rect 720 950 724 970
rect 728 950 732 970
rect 736 950 740 970
rect 797 950 801 970
rect 805 950 809 970
rect 813 950 817 970
rect 862 950 866 970
rect 870 950 874 970
rect 878 950 882 970
rect 937 950 941 970
rect 945 950 949 970
rect 953 950 957 970
rect 1002 950 1006 970
rect 1010 950 1014 970
rect 1018 950 1022 970
rect 1082 950 1086 970
rect 1090 950 1094 970
rect 1098 950 1102 970
rect 1147 950 1151 970
rect 1155 950 1159 970
rect 1163 950 1167 970
rect 1227 950 1231 970
rect 1235 950 1239 970
rect 1243 950 1247 970
rect 1292 950 1296 970
rect 1300 950 1304 970
rect 1308 950 1312 970
rect 1372 950 1376 970
rect 1380 950 1384 970
rect 1388 950 1392 970
rect 1437 950 1441 970
rect 1445 950 1449 970
rect 1453 950 1457 970
rect -248 940 -228 944
rect -575 932 -555 936
rect 165 940 185 944
rect -248 932 -228 936
rect 165 932 185 936
rect 165 924 185 928
rect -1330 904 -1326 924
rect -1322 904 -1318 924
rect -1279 904 -1275 924
rect -1271 904 -1267 924
rect -1234 905 -1214 909
rect -1128 905 -1108 909
rect -1234 897 -1214 901
rect -1002 904 -998 924
rect -994 904 -990 924
rect -952 904 -948 924
rect -944 904 -940 924
rect -907 905 -887 909
rect -1128 897 -1108 901
rect -1234 889 -1214 893
rect -1128 889 -1108 893
rect -801 905 -781 909
rect -907 897 -887 901
rect -801 897 -781 901
rect -907 889 -887 893
rect -671 900 -667 920
rect -663 900 -659 920
rect -620 900 -616 920
rect -612 900 -608 920
rect -575 901 -555 905
rect -801 889 -781 893
rect -469 901 -449 905
rect -575 893 -555 897
rect -343 900 -339 920
rect -335 900 -331 920
rect -293 900 -289 920
rect -285 900 -281 920
rect 74 906 94 910
rect -248 901 -228 905
rect -469 893 -449 897
rect -575 885 -555 889
rect -469 885 -449 889
rect -142 901 -122 905
rect -248 893 -228 897
rect 261 906 281 910
rect 74 898 94 902
rect -142 893 -122 897
rect -248 885 -228 889
rect 261 898 281 902
rect 74 890 94 894
rect 261 890 281 894
rect 441 892 445 912
rect 449 892 453 912
rect 569 892 573 912
rect 577 892 581 912
rect -142 885 -122 889
rect 165 884 185 888
rect 368 887 388 891
rect 165 876 185 880
rect 368 879 388 883
rect 486 886 526 890
rect 486 878 526 882
rect 165 868 185 872
rect 368 871 388 875
rect 486 870 526 874
rect 132 831 136 851
rect 140 831 144 851
rect 673 844 677 864
rect 681 844 685 864
rect 689 844 693 864
rect 720 844 724 864
rect 728 844 732 864
rect 736 844 740 864
rect 815 844 819 864
rect 823 844 827 864
rect 831 844 835 864
rect 862 844 866 864
rect 870 844 874 864
rect 878 844 882 864
rect 955 844 959 864
rect 963 844 967 864
rect 971 844 975 864
rect 1002 844 1006 864
rect 1010 844 1014 864
rect 1018 844 1022 864
rect 1100 844 1104 864
rect 1108 844 1112 864
rect 1116 844 1120 864
rect 1147 844 1151 864
rect 1155 844 1159 864
rect 1163 844 1167 864
rect 1245 844 1249 864
rect 1253 844 1257 864
rect 1261 844 1265 864
rect 1292 844 1296 864
rect 1300 844 1304 864
rect 1308 844 1312 864
rect 1390 844 1394 864
rect 1398 844 1402 864
rect 1406 844 1410 864
rect 1437 844 1441 864
rect 1445 844 1449 864
rect 1453 844 1457 864
rect 59 826 79 830
rect 59 818 79 822
rect 59 810 79 814
rect 364 806 368 826
rect 372 806 376 826
rect 291 801 311 805
rect 291 793 311 797
rect 415 804 475 808
rect 415 796 475 800
rect 517 799 521 819
rect 525 799 529 819
rect 705 807 725 811
rect 847 807 867 811
rect 987 807 1007 811
rect 1132 807 1152 811
rect 1277 807 1297 811
rect 1422 807 1442 811
rect 705 799 725 803
rect 847 799 867 803
rect 987 799 1007 803
rect 1132 799 1152 803
rect 1277 799 1297 803
rect 1422 799 1442 803
rect 291 785 311 789
rect 415 788 475 792
rect 415 780 475 784
rect 164 760 184 764
rect 164 752 184 756
rect 705 756 725 760
rect 847 756 867 760
rect 987 756 1007 760
rect 1132 756 1152 760
rect 1277 756 1297 760
rect 1422 756 1442 760
rect 164 744 184 748
rect 705 748 725 752
rect 847 748 867 752
rect 987 748 1007 752
rect 1132 748 1152 752
rect 1277 748 1297 752
rect 1422 748 1442 752
rect -1128 731 -1108 735
rect -801 731 -781 735
rect -1128 723 -1108 727
rect -469 730 -449 734
rect -801 723 -781 727
rect -1234 713 -1214 717
rect -1128 715 -1108 719
rect -142 730 -122 734
rect -469 722 -449 726
rect -907 713 -887 717
rect -1234 705 -1214 709
rect -801 715 -781 719
rect -142 722 -122 726
rect -575 712 -555 716
rect -907 705 -887 709
rect -1234 697 -1214 701
rect -469 714 -449 718
rect 73 726 93 730
rect 260 726 280 730
rect -248 712 -228 716
rect -575 704 -555 708
rect -907 697 -887 701
rect -142 714 -122 718
rect 73 718 93 722
rect 260 718 280 722
rect 73 710 93 714
rect 374 719 394 723
rect 260 710 280 714
rect 374 711 394 715
rect -248 704 -228 708
rect -575 696 -555 700
rect 164 704 184 708
rect -248 696 -228 700
rect 456 713 460 733
rect 464 713 468 733
rect 374 703 394 707
rect 164 696 184 700
rect 374 695 394 699
rect 164 688 184 692
rect -1330 665 -1326 685
rect -1322 665 -1318 685
rect -1279 665 -1275 685
rect -1271 665 -1267 685
rect -1234 666 -1214 670
rect -1128 666 -1108 670
rect -1234 658 -1214 662
rect -1002 665 -998 685
rect -994 665 -990 685
rect -952 665 -948 685
rect -944 665 -940 685
rect -907 666 -887 670
rect -1128 658 -1108 662
rect -1234 650 -1214 654
rect -1128 650 -1108 654
rect -801 666 -781 670
rect -907 658 -887 662
rect -671 664 -667 684
rect -663 664 -659 684
rect -620 664 -616 684
rect -612 664 -608 684
rect -575 665 -555 669
rect -801 658 -781 662
rect -907 650 -887 654
rect -801 650 -781 654
rect -469 665 -449 669
rect -575 657 -555 661
rect -343 664 -339 684
rect -335 664 -331 684
rect -293 664 -289 684
rect -285 664 -281 684
rect 655 673 675 677
rect -248 665 -228 669
rect -469 657 -449 661
rect -575 649 -555 653
rect -469 649 -449 653
rect -142 665 -122 669
rect -248 657 -228 661
rect -142 657 -122 661
rect -248 649 -228 653
rect -142 649 -122 653
rect 131 651 135 671
rect 139 651 143 671
rect 655 665 675 669
rect 655 657 675 661
rect 58 646 78 650
rect 58 638 78 642
rect 564 639 584 643
rect 58 630 78 634
rect 296 633 316 637
rect 751 639 771 643
rect 564 631 584 635
rect 296 625 316 629
rect 751 631 771 635
rect 564 623 584 627
rect 751 623 771 627
rect 296 617 316 621
rect 655 617 675 621
rect 655 609 675 613
rect 205 599 225 603
rect 392 599 412 603
rect 205 591 225 595
rect 655 601 675 605
rect 392 591 412 595
rect 205 583 225 587
rect 392 583 412 587
rect 296 577 316 581
rect 296 569 316 573
rect 296 561 316 565
rect 621 540 625 560
rect 629 540 633 560
rect 548 535 568 539
rect 548 527 568 531
rect -1128 517 -1108 521
rect -801 517 -781 521
rect -1128 509 -1108 513
rect -469 516 -449 520
rect -801 509 -781 513
rect -1234 499 -1214 503
rect -1128 501 -1108 505
rect -142 516 -122 520
rect -469 508 -449 512
rect -907 499 -887 503
rect -1234 491 -1214 495
rect -801 501 -781 505
rect 548 519 568 523
rect -142 508 -122 512
rect -575 498 -555 502
rect -907 491 -887 495
rect -1234 483 -1214 487
rect -469 500 -449 504
rect 164 506 184 510
rect -248 498 -228 502
rect -575 490 -555 494
rect -907 483 -887 487
rect -142 500 -122 504
rect 164 498 184 502
rect -248 490 -228 494
rect -575 482 -555 486
rect 695 498 775 502
rect 164 490 184 494
rect -248 482 -228 486
rect 379 484 399 488
rect 379 476 399 480
rect -1330 451 -1326 471
rect -1322 451 -1318 471
rect -1279 451 -1275 471
rect -1271 451 -1267 471
rect -1234 452 -1214 456
rect -1128 452 -1108 456
rect -1234 444 -1214 448
rect -1002 451 -998 471
rect -994 451 -990 471
rect -952 451 -948 471
rect -944 451 -940 471
rect 73 472 93 476
rect -907 452 -887 456
rect -1128 444 -1108 448
rect -1234 436 -1214 440
rect -1128 436 -1108 440
rect -801 452 -781 456
rect -907 444 -887 448
rect -671 450 -667 470
rect -663 450 -659 470
rect -620 450 -616 470
rect -612 450 -608 470
rect -575 451 -555 455
rect -801 444 -781 448
rect -907 436 -887 440
rect -801 436 -781 440
rect -469 451 -449 455
rect -575 443 -555 447
rect -343 450 -339 470
rect -335 450 -331 470
rect -293 450 -289 470
rect -285 450 -281 470
rect 260 472 280 476
rect 73 464 93 468
rect 471 475 475 495
rect 479 475 483 495
rect 548 482 568 486
rect 260 464 280 468
rect 73 456 93 460
rect 379 468 399 472
rect 260 456 280 460
rect 379 460 399 464
rect 548 474 568 478
rect 630 476 634 496
rect 638 476 642 496
rect 695 490 775 494
rect 818 487 822 507
rect 826 487 830 507
rect 695 482 775 486
rect 548 466 568 470
rect -248 451 -228 455
rect -469 443 -449 447
rect -575 435 -555 439
rect -469 435 -449 439
rect -142 451 -122 455
rect -248 443 -228 447
rect 164 450 184 454
rect -142 443 -122 447
rect -248 435 -228 439
rect 379 452 399 456
rect 548 458 568 462
rect 695 474 775 478
rect 695 466 775 470
rect 164 442 184 446
rect -142 435 -122 439
rect 164 434 184 438
rect 798 419 802 439
rect 806 419 810 439
rect 131 397 135 417
rect 139 397 143 417
rect 725 414 745 418
rect 725 406 745 410
rect 725 398 745 402
rect 58 392 78 396
rect 58 384 78 388
rect 58 376 78 380
rect 307 371 327 375
rect 307 363 327 367
rect 385 363 389 383
rect 393 363 397 383
rect 443 373 463 377
rect 443 365 463 369
rect 307 355 327 359
rect 307 347 327 351
rect 535 364 539 384
rect 543 364 547 384
rect 589 370 609 374
rect 443 357 463 361
rect 443 349 463 353
rect 307 339 327 343
rect 589 362 609 366
rect 671 364 675 384
rect 679 364 683 384
rect 589 354 609 358
rect 443 341 463 345
rect 589 346 609 350
rect 735 350 835 354
rect 735 342 835 346
rect 876 343 880 363
rect 884 343 888 363
rect 307 331 327 335
rect 735 334 835 338
rect 165 324 185 328
rect 735 326 835 330
rect 165 316 185 320
rect 735 318 835 322
rect 165 308 185 312
rect 735 310 835 314
rect 74 290 94 294
rect 261 290 281 294
rect 74 282 94 286
rect -1128 278 -1108 282
rect -801 278 -781 282
rect -1128 270 -1108 274
rect -469 277 -449 281
rect -801 270 -781 274
rect -1234 260 -1214 264
rect -1128 262 -1108 266
rect -142 277 -122 281
rect -469 269 -449 273
rect -907 260 -887 264
rect -1234 252 -1214 256
rect -801 262 -781 266
rect 261 282 281 286
rect 74 274 94 278
rect 261 274 281 278
rect -142 269 -122 273
rect -575 259 -555 263
rect -907 252 -887 256
rect -1234 244 -1214 248
rect -469 261 -449 265
rect 165 268 185 272
rect -248 259 -228 263
rect -575 251 -555 255
rect -907 244 -887 248
rect -142 261 -122 265
rect 165 260 185 264
rect -248 251 -228 255
rect -575 243 -555 247
rect 165 252 185 256
rect 488 255 508 259
rect 1113 252 1133 256
rect -248 243 -228 247
rect 488 247 508 251
rect 1113 244 1133 248
rect 488 239 508 243
rect -1330 212 -1326 232
rect -1322 212 -1318 232
rect -1279 212 -1275 232
rect -1271 212 -1267 232
rect -1234 213 -1214 217
rect -1128 213 -1108 217
rect -1234 205 -1214 209
rect -1002 212 -998 232
rect -994 212 -990 232
rect -952 212 -948 232
rect -944 212 -940 232
rect -907 213 -887 217
rect -1128 205 -1108 209
rect -1234 197 -1214 201
rect -1128 197 -1108 201
rect -801 213 -781 217
rect -907 205 -887 209
rect -671 211 -667 231
rect -663 211 -659 231
rect -620 211 -616 231
rect -612 211 -608 231
rect -575 212 -555 216
rect -801 205 -781 209
rect -907 197 -887 201
rect -801 197 -781 201
rect -469 212 -449 216
rect -575 204 -555 208
rect -343 211 -339 231
rect -335 211 -331 231
rect -293 211 -289 231
rect -285 211 -281 231
rect -248 212 -228 216
rect -469 204 -449 208
rect -575 196 -555 200
rect -469 196 -449 200
rect -142 212 -122 216
rect -248 204 -228 208
rect 132 215 136 235
rect 140 215 144 235
rect 397 221 417 225
rect 584 221 604 225
rect 59 210 79 214
rect -142 204 -122 208
rect -248 196 -228 200
rect 59 202 79 206
rect -142 196 -122 200
rect 397 213 417 217
rect 925 219 929 239
rect 933 219 937 239
rect 1113 236 1133 240
rect 584 213 604 217
rect 397 205 417 209
rect 584 205 604 209
rect 488 199 508 203
rect 59 194 79 198
rect 706 202 726 206
rect 488 191 508 195
rect 706 194 726 198
rect 788 196 792 216
rect 796 196 800 216
rect 852 214 872 218
rect 852 206 872 210
rect 1022 218 1042 222
rect 1209 218 1229 222
rect 1022 210 1042 214
rect 1209 210 1229 214
rect 852 198 872 202
rect 488 183 508 187
rect 706 186 726 190
rect 706 178 726 182
rect 1022 202 1042 206
rect 1209 202 1229 206
rect 1113 196 1133 200
rect 1113 188 1133 192
rect 1113 180 1133 184
rect 166 141 186 145
rect 166 133 186 137
rect 389 131 399 135
rect 166 125 186 129
rect 389 123 399 127
rect 389 115 399 119
rect 470 116 474 136
rect 478 116 482 136
rect 525 133 545 137
rect 525 125 545 129
rect 603 125 607 145
rect 611 125 615 145
rect 653 125 673 129
rect 525 117 545 121
rect 75 107 95 111
rect 262 107 282 111
rect 75 99 95 103
rect 389 107 399 111
rect 262 99 282 103
rect -1128 91 -1108 95
rect -801 91 -781 95
rect -1128 83 -1108 87
rect -469 90 -449 94
rect -801 83 -781 87
rect -1234 73 -1214 77
rect -1128 75 -1108 79
rect -142 90 -122 94
rect -469 82 -449 86
rect -907 73 -887 77
rect -1234 65 -1214 69
rect -801 75 -781 79
rect 75 91 95 95
rect 389 99 399 103
rect 262 91 282 95
rect 525 109 545 113
rect 653 117 673 121
rect 745 116 749 136
rect 753 116 757 136
rect 864 129 984 133
rect 864 121 984 125
rect 653 109 673 113
rect 525 101 545 105
rect 389 91 399 95
rect -142 82 -122 86
rect -575 72 -555 76
rect -907 65 -887 69
rect -1234 57 -1214 61
rect -469 74 -449 78
rect 166 85 186 89
rect 653 101 673 105
rect 525 93 545 97
rect 864 113 984 117
rect 1034 114 1038 134
rect 1042 114 1046 134
rect 864 105 984 109
rect 653 93 673 97
rect 864 97 984 101
rect 389 83 399 87
rect 864 89 984 93
rect -248 72 -228 76
rect -575 64 -555 68
rect -907 57 -887 61
rect -142 74 -122 78
rect 166 77 186 81
rect 864 81 984 85
rect 166 69 186 73
rect -248 64 -228 68
rect -575 56 -555 60
rect -248 56 -228 60
rect -1330 25 -1326 45
rect -1322 25 -1318 45
rect -1279 25 -1275 45
rect -1271 25 -1267 45
rect -1234 26 -1214 30
rect -1128 26 -1108 30
rect -1234 18 -1214 22
rect -1002 25 -998 45
rect -994 25 -990 45
rect -952 25 -948 45
rect -944 25 -940 45
rect -907 26 -887 30
rect -1128 18 -1108 22
rect -1234 10 -1214 14
rect -1128 10 -1108 14
rect -801 26 -781 30
rect -907 18 -887 22
rect -671 24 -667 44
rect -663 24 -659 44
rect -620 24 -616 44
rect -612 24 -608 44
rect -575 25 -555 29
rect -801 18 -781 22
rect -907 10 -887 14
rect -801 10 -781 14
rect -469 25 -449 29
rect -575 17 -555 21
rect -343 24 -339 44
rect -335 24 -331 44
rect -293 24 -289 44
rect -285 24 -281 44
rect 133 32 137 52
rect 141 32 145 52
rect -248 25 -228 29
rect -469 17 -449 21
rect -575 9 -555 13
rect -469 9 -449 13
rect -142 25 -122 29
rect -248 17 -228 21
rect 60 27 80 31
rect -142 17 -122 21
rect -248 9 -228 13
rect 60 19 80 23
rect -142 9 -122 13
rect 60 11 80 15
<< m2contact >>
rect 654 1352 659 1357
rect 654 1335 659 1340
rect 678 1304 683 1310
rect 693 1304 698 1310
rect 709 1268 714 1273
rect 644 1251 649 1256
rect 678 1259 683 1264
rect 695 1232 700 1237
rect 713 1233 718 1238
rect 796 1352 801 1357
rect 796 1335 801 1340
rect 820 1304 825 1310
rect -494 1140 -489 1145
rect -646 1099 -641 1104
rect -656 1090 -651 1095
rect -599 1099 -594 1104
rect -625 1090 -620 1095
rect -606 1090 -601 1095
rect -410 1130 -405 1135
rect -486 1106 -481 1111
rect -441 1106 -435 1111
rect -393 1130 -388 1135
rect -585 1088 -580 1093
rect -513 1089 -508 1094
rect -585 1072 -580 1077
rect -512 1071 -507 1076
rect -441 1091 -435 1096
rect -477 1075 -472 1080
rect -261 1122 -256 1128
rect -167 1140 -162 1145
rect -318 1099 -313 1104
rect -336 1094 -331 1099
rect -358 1052 -353 1057
rect -272 1099 -267 1104
rect -298 1090 -293 1095
rect -279 1090 -274 1095
rect -83 1130 -78 1135
rect -159 1106 -154 1111
rect -114 1106 -108 1111
rect -66 1130 -61 1135
rect -258 1088 -253 1093
rect -186 1089 -181 1094
rect -258 1072 -253 1077
rect -185 1071 -180 1076
rect -114 1091 -108 1096
rect -150 1075 -145 1080
rect -1154 980 -1149 985
rect -1306 939 -1301 944
rect -1316 930 -1311 935
rect -1259 939 -1254 944
rect -1285 930 -1280 935
rect -1266 930 -1261 935
rect -1070 970 -1065 975
rect -1146 946 -1141 951
rect -1101 946 -1095 951
rect -1053 970 -1048 975
rect -1245 928 -1240 933
rect -1173 929 -1168 934
rect -1245 912 -1240 917
rect -1172 911 -1167 916
rect -1101 931 -1095 936
rect -1137 915 -1132 920
rect -921 962 -916 968
rect -827 980 -822 985
rect -978 939 -973 944
rect -996 934 -991 939
rect -1018 892 -1013 897
rect -932 939 -927 944
rect -958 930 -953 935
rect -939 930 -934 935
rect -743 970 -738 975
rect -819 946 -814 951
rect -774 946 -768 951
rect -726 970 -721 975
rect -918 928 -913 933
rect -846 929 -841 934
rect -918 912 -913 917
rect -845 911 -840 916
rect -774 931 -768 936
rect -810 915 -805 920
rect -495 976 -490 981
rect -647 935 -642 940
rect -657 926 -652 931
rect -600 935 -595 940
rect -626 926 -621 931
rect -607 926 -602 931
rect -411 966 -406 971
rect -487 942 -482 947
rect -442 942 -436 947
rect -394 966 -389 971
rect -586 924 -581 929
rect -514 925 -509 930
rect -586 908 -581 913
rect -513 907 -508 912
rect -442 927 -436 932
rect -478 911 -473 916
rect -262 958 -257 964
rect -168 976 -163 981
rect -319 935 -314 940
rect -337 930 -332 935
rect -359 888 -354 893
rect -273 935 -268 940
rect -299 926 -294 931
rect -280 926 -275 931
rect -84 966 -79 971
rect -160 942 -155 947
rect -115 942 -109 947
rect -67 966 -62 971
rect -259 924 -254 929
rect -187 925 -182 930
rect -259 908 -254 913
rect -186 907 -181 912
rect -115 927 -109 932
rect -151 911 -146 916
rect 315 1041 320 1046
rect 475 1027 480 1032
rect 315 998 320 1003
rect 64 953 69 958
rect 224 939 229 944
rect 64 910 69 915
rect 14 894 19 899
rect 42 894 47 899
rect 134 905 139 910
rect 205 911 210 916
rect 385 993 390 998
rect 289 963 294 968
rect 456 999 461 1004
rect 501 998 506 1003
rect 572 994 577 999
rect 335 920 340 925
rect 250 910 255 915
rect 321 906 326 911
rect 344 892 349 897
rect 334 865 340 871
rect 23 818 28 823
rect 446 846 451 851
rect 63 773 68 778
rect -1154 741 -1149 746
rect -1306 700 -1301 705
rect -1316 691 -1311 696
rect -1259 700 -1254 705
rect -1285 691 -1280 696
rect -1266 691 -1261 696
rect -1070 731 -1065 736
rect -1146 707 -1141 712
rect -1101 707 -1095 712
rect -1053 731 -1048 736
rect -1245 689 -1240 694
rect -1173 690 -1168 695
rect -1245 673 -1240 678
rect -1172 672 -1167 677
rect -1101 692 -1095 697
rect -1137 676 -1132 681
rect -921 723 -916 729
rect -827 741 -822 746
rect -978 700 -973 705
rect -996 695 -991 700
rect -1018 653 -1013 658
rect -932 700 -927 705
rect -958 691 -953 696
rect -939 691 -934 696
rect -743 731 -738 736
rect -819 707 -814 712
rect -774 707 -768 712
rect -726 731 -721 736
rect -918 689 -913 694
rect -846 690 -841 695
rect -918 673 -913 678
rect -845 672 -840 677
rect -774 692 -768 697
rect -810 676 -805 681
rect -495 740 -490 745
rect -647 699 -642 704
rect -657 690 -652 695
rect -600 699 -595 704
rect -626 690 -621 695
rect -607 690 -602 695
rect -411 730 -406 735
rect -487 706 -482 711
rect -442 706 -436 711
rect -394 730 -389 735
rect -586 688 -581 693
rect -514 689 -509 694
rect -586 672 -581 677
rect -513 671 -508 676
rect -442 691 -436 696
rect -478 675 -473 680
rect -262 722 -257 728
rect -168 740 -163 745
rect -319 699 -314 704
rect -337 694 -332 699
rect -359 652 -354 657
rect -273 699 -268 704
rect -299 690 -294 695
rect -280 690 -275 695
rect -84 730 -79 735
rect -160 706 -155 711
rect -115 706 -109 711
rect -67 730 -62 735
rect -259 688 -254 693
rect -187 689 -182 694
rect -259 672 -254 677
rect -186 671 -181 676
rect -115 691 -109 696
rect -151 675 -146 680
rect 223 759 228 764
rect 63 730 68 735
rect 13 714 18 719
rect 41 714 46 719
rect 133 725 138 730
rect 204 731 209 736
rect 533 786 538 791
rect 249 730 254 735
rect 320 726 325 731
rect 288 692 293 697
rect 330 712 335 717
rect 344 698 349 703
rect 439 702 444 707
rect 22 638 27 643
rect 195 646 200 651
rect 167 599 172 604
rect 355 632 360 637
rect 195 603 200 608
rect 265 598 270 603
rect -1154 527 -1149 532
rect -1306 486 -1301 491
rect -1316 477 -1311 482
rect -1259 486 -1254 491
rect -1285 477 -1280 482
rect -1266 477 -1261 482
rect -1070 517 -1065 522
rect -1146 493 -1141 498
rect -1101 493 -1095 498
rect -1053 517 -1048 522
rect -1245 475 -1240 480
rect -1173 476 -1168 481
rect -1245 459 -1240 464
rect -1172 458 -1167 463
rect -1101 478 -1095 483
rect -1137 462 -1132 467
rect -921 509 -916 515
rect -827 527 -822 532
rect -978 486 -973 491
rect -996 481 -991 486
rect -1018 439 -1013 444
rect -932 486 -927 491
rect -958 477 -953 482
rect -939 477 -934 482
rect -743 517 -738 522
rect -819 493 -814 498
rect -774 493 -768 498
rect -726 517 -721 522
rect -918 475 -913 480
rect -846 476 -841 481
rect -918 459 -913 464
rect -845 458 -840 463
rect -774 478 -768 483
rect -810 462 -805 467
rect -495 526 -490 531
rect -647 485 -642 490
rect -657 476 -652 481
rect -600 485 -595 490
rect -626 476 -621 481
rect -607 476 -602 481
rect -411 516 -406 521
rect -487 492 -482 497
rect -442 492 -436 497
rect -394 516 -389 521
rect -586 474 -581 479
rect -514 475 -509 480
rect -586 458 -581 463
rect -513 457 -508 462
rect -442 477 -436 482
rect -478 461 -473 466
rect -262 508 -257 514
rect -168 526 -163 531
rect -319 485 -314 490
rect -337 480 -332 485
rect -359 438 -354 443
rect -273 485 -268 490
rect -299 476 -294 481
rect -280 476 -275 481
rect -84 516 -79 521
rect -160 492 -155 497
rect -115 492 -109 497
rect -67 516 -62 521
rect -259 474 -254 479
rect -187 475 -182 480
rect -259 458 -254 463
rect -186 457 -181 462
rect -115 477 -109 482
rect -151 461 -146 466
rect 336 604 341 609
rect 381 603 386 608
rect 452 599 457 604
rect 489 559 494 564
rect 470 552 475 557
rect 661 1157 667 1162
rect 696 1160 701 1165
rect 712 1160 717 1165
rect 685 1146 690 1151
rect 694 1139 699 1144
rect 835 1304 840 1310
rect 851 1268 856 1273
rect 786 1251 791 1256
rect 820 1259 825 1264
rect 837 1232 842 1237
rect 855 1233 860 1238
rect 936 1352 941 1357
rect 936 1335 941 1340
rect 960 1304 965 1310
rect 694 1120 699 1125
rect 685 1100 690 1105
rect 690 1082 695 1087
rect 732 1060 737 1065
rect 654 1025 659 1030
rect 654 1008 659 1013
rect 678 977 683 983
rect 693 977 698 983
rect 709 941 714 946
rect 644 924 649 929
rect 678 932 683 937
rect 695 905 700 910
rect 713 906 718 911
rect 696 833 701 838
rect 712 833 717 838
rect 685 819 690 824
rect 694 812 699 817
rect 803 1157 809 1162
rect 838 1160 843 1165
rect 854 1160 859 1165
rect 827 1146 832 1151
rect 836 1139 841 1144
rect 975 1304 980 1310
rect 991 1268 996 1273
rect 926 1251 931 1256
rect 960 1259 965 1264
rect 977 1232 982 1237
rect 995 1233 1000 1238
rect 1081 1352 1086 1357
rect 1081 1335 1086 1340
rect 1105 1304 1110 1310
rect 836 1120 841 1125
rect 827 1100 832 1105
rect 832 1082 837 1087
rect 874 1060 879 1065
rect 796 1025 801 1030
rect 796 1008 801 1013
rect 820 977 825 983
rect 835 977 840 983
rect 851 941 856 946
rect 786 924 791 929
rect 694 793 699 798
rect 685 772 690 777
rect 694 762 699 767
rect 820 932 825 937
rect 837 905 842 910
rect 855 906 860 911
rect 838 833 843 838
rect 854 833 859 838
rect 827 819 832 824
rect 836 812 841 817
rect 943 1157 949 1162
rect 978 1160 983 1165
rect 994 1160 999 1165
rect 967 1146 972 1151
rect 976 1139 981 1144
rect 1120 1304 1125 1310
rect 1136 1268 1141 1273
rect 1071 1251 1076 1256
rect 1105 1259 1110 1264
rect 1122 1232 1127 1237
rect 1140 1233 1145 1238
rect 1226 1352 1231 1357
rect 1226 1335 1231 1340
rect 1250 1304 1255 1310
rect 976 1120 981 1125
rect 967 1100 972 1105
rect 972 1082 977 1087
rect 1014 1060 1019 1065
rect 936 1025 941 1030
rect 936 1008 941 1013
rect 960 977 965 983
rect 975 977 980 983
rect 991 941 996 946
rect 926 924 931 929
rect 836 793 841 798
rect 827 772 832 777
rect 836 762 841 767
rect 819 728 824 733
rect 960 932 965 937
rect 977 905 982 910
rect 995 906 1000 911
rect 978 833 983 838
rect 994 833 999 838
rect 967 819 972 824
rect 976 812 981 817
rect 1088 1157 1094 1162
rect 1123 1160 1128 1165
rect 1139 1160 1144 1165
rect 1112 1146 1117 1151
rect 1121 1139 1126 1144
rect 1265 1304 1270 1310
rect 1281 1268 1286 1273
rect 1216 1251 1221 1256
rect 1250 1259 1255 1264
rect 1267 1232 1272 1237
rect 1285 1233 1290 1238
rect 1371 1352 1376 1357
rect 1371 1335 1376 1340
rect 1395 1304 1400 1310
rect 1121 1120 1126 1125
rect 1112 1100 1117 1105
rect 1117 1082 1122 1087
rect 1159 1060 1164 1065
rect 1081 1025 1086 1030
rect 1081 1008 1086 1013
rect 1105 977 1110 983
rect 1120 977 1125 983
rect 1136 941 1141 946
rect 1071 924 1076 929
rect 976 793 981 798
rect 554 686 559 691
rect 531 636 536 641
rect 714 672 719 677
rect 554 643 559 648
rect 624 638 629 643
rect 63 519 68 524
rect 223 505 228 510
rect 63 476 68 481
rect 13 460 18 465
rect 41 460 46 465
rect 133 471 138 476
rect 204 477 209 482
rect 369 530 374 535
rect 470 531 475 536
rect 695 644 700 649
rect 740 643 745 648
rect 967 772 972 777
rect 976 762 981 767
rect 1105 932 1110 937
rect 1122 905 1127 910
rect 1140 906 1145 911
rect 1123 833 1128 838
rect 1139 833 1144 838
rect 1112 819 1117 824
rect 1121 812 1126 817
rect 1233 1157 1239 1162
rect 1268 1160 1273 1165
rect 1284 1160 1289 1165
rect 1257 1146 1262 1151
rect 1266 1139 1271 1144
rect 1410 1304 1415 1310
rect 1426 1268 1431 1273
rect 1361 1251 1366 1256
rect 1395 1259 1400 1264
rect 1412 1232 1417 1237
rect 1430 1233 1435 1238
rect 1266 1120 1271 1125
rect 1257 1100 1262 1105
rect 1262 1082 1267 1087
rect 1304 1060 1309 1065
rect 1226 1025 1231 1030
rect 1226 1008 1231 1013
rect 1250 977 1255 983
rect 1265 977 1270 983
rect 1281 941 1286 946
rect 1216 924 1221 929
rect 1121 793 1126 798
rect 1112 772 1117 777
rect 1121 762 1126 767
rect 1250 932 1255 937
rect 1267 905 1272 910
rect 1285 906 1290 911
rect 1268 833 1273 838
rect 1284 833 1289 838
rect 1257 819 1262 824
rect 1266 812 1271 817
rect 1378 1157 1384 1162
rect 1413 1160 1418 1165
rect 1429 1160 1434 1165
rect 1402 1146 1407 1151
rect 1411 1139 1416 1144
rect 1411 1120 1416 1125
rect 1402 1100 1407 1105
rect 1407 1082 1412 1087
rect 1449 1060 1454 1065
rect 1371 1025 1376 1030
rect 1371 1008 1376 1013
rect 1395 977 1400 983
rect 1410 977 1415 983
rect 1426 941 1431 946
rect 1361 924 1366 929
rect 1266 793 1271 798
rect 811 639 816 644
rect 1257 772 1262 777
rect 1266 762 1271 767
rect 1395 932 1400 937
rect 1412 905 1417 910
rect 1430 906 1435 911
rect 1413 833 1418 838
rect 1429 833 1434 838
rect 1402 819 1407 824
rect 1411 812 1416 817
rect 1411 793 1416 798
rect 1402 772 1407 777
rect 1411 762 1416 767
rect 531 545 536 550
rect 496 517 501 522
rect 341 507 346 512
rect 350 491 355 496
rect 362 488 367 493
rect 249 476 254 481
rect 341 481 346 486
rect 320 472 325 477
rect 354 475 359 480
rect 341 465 346 470
rect 501 483 506 488
rect 522 487 527 492
rect 454 459 459 464
rect 512 471 517 476
rect 655 485 661 491
rect 493 441 499 447
rect 506 446 511 451
rect 331 431 336 436
rect 22 384 27 389
rect 506 405 511 410
rect 695 402 700 407
rect 781 405 787 411
rect 853 455 858 460
rect 853 427 858 432
rect 838 413 843 418
rect 289 379 294 384
rect 278 369 283 374
rect 268 358 273 363
rect 259 347 264 352
rect 64 337 69 342
rect -1154 288 -1149 293
rect -1306 247 -1301 252
rect -1316 238 -1311 243
rect -1259 247 -1254 252
rect -1285 238 -1280 243
rect -1266 238 -1261 243
rect -1070 278 -1065 283
rect -1146 254 -1141 259
rect -1101 254 -1095 259
rect -1053 278 -1048 283
rect -1245 236 -1240 241
rect -1173 237 -1168 242
rect -1245 220 -1240 225
rect -1172 219 -1167 224
rect -1101 239 -1095 244
rect -1137 223 -1132 228
rect -921 270 -916 276
rect -827 288 -822 293
rect -978 247 -973 252
rect -996 242 -991 247
rect -1018 200 -1013 205
rect -932 247 -927 252
rect -958 238 -953 243
rect -939 238 -934 243
rect -743 278 -738 283
rect -819 254 -814 259
rect -774 254 -768 259
rect -726 278 -721 283
rect -918 236 -913 241
rect -846 237 -841 242
rect -918 220 -913 225
rect -845 219 -840 224
rect -774 239 -768 244
rect -810 223 -805 228
rect -495 287 -490 292
rect -647 246 -642 251
rect -657 237 -652 242
rect -600 246 -595 251
rect -626 237 -621 242
rect -607 237 -602 242
rect -411 277 -406 282
rect -487 253 -482 258
rect -442 253 -436 258
rect -394 277 -389 282
rect -586 235 -581 240
rect -514 236 -509 241
rect -586 219 -581 224
rect -513 218 -508 223
rect -442 238 -436 243
rect -478 222 -473 227
rect -262 269 -257 275
rect -168 287 -163 292
rect -319 246 -314 251
rect -337 241 -332 246
rect -359 199 -354 204
rect -273 246 -268 251
rect -299 237 -294 242
rect -280 237 -275 242
rect -84 277 -79 282
rect -160 253 -155 258
rect -115 253 -109 258
rect 224 323 229 328
rect 64 294 69 299
rect -67 277 -62 282
rect 14 278 19 283
rect -259 235 -254 240
rect -187 236 -182 241
rect -259 219 -254 224
rect -186 218 -181 223
rect -115 238 -109 243
rect -151 222 -146 227
rect 42 278 47 283
rect 134 289 139 294
rect 205 295 210 300
rect 422 377 427 382
rect 404 359 409 364
rect 367 346 372 351
rect 269 305 275 311
rect 375 332 380 337
rect 413 349 418 354
rect 563 376 568 381
rect 554 358 559 363
rect 518 348 523 353
rect 425 332 430 337
rect 654 354 659 359
rect 826 400 831 405
rect 894 386 899 391
rect 697 374 702 379
rect 819 372 824 377
rect 688 351 693 356
rect 569 336 574 341
rect 706 338 711 343
rect 705 329 710 334
rect 366 313 371 318
rect 461 315 466 320
rect 556 315 562 321
rect 250 294 255 299
rect 321 290 326 295
rect 256 258 262 264
rect 288 258 294 264
rect 387 268 392 273
rect 23 202 28 207
rect 257 229 262 234
rect 269 227 275 233
rect 311 224 317 230
rect 547 254 552 259
rect 387 225 392 230
rect 336 214 341 219
rect 457 220 462 225
rect 280 199 285 204
rect 65 154 70 159
rect -1154 101 -1149 106
rect -1306 60 -1301 65
rect -1316 51 -1311 56
rect -1259 60 -1254 65
rect -1285 51 -1280 56
rect -1266 51 -1261 56
rect -1070 91 -1065 96
rect -1146 67 -1141 72
rect -1101 67 -1095 72
rect -1053 91 -1048 96
rect -1245 49 -1240 54
rect -1173 50 -1168 55
rect -1245 33 -1240 38
rect -1172 32 -1167 37
rect -1101 52 -1095 57
rect -1137 36 -1132 41
rect -921 83 -916 89
rect -827 101 -822 106
rect -978 60 -973 65
rect -996 55 -991 60
rect -1018 13 -1013 18
rect -932 60 -927 65
rect -958 51 -953 56
rect -939 51 -934 56
rect -743 91 -738 96
rect -819 67 -814 72
rect -774 67 -768 72
rect -726 91 -721 96
rect -918 49 -913 54
rect -846 50 -841 55
rect -918 33 -913 38
rect -845 32 -840 37
rect -774 52 -768 57
rect -810 36 -805 41
rect -495 100 -490 105
rect -647 59 -642 64
rect -657 50 -652 55
rect -600 59 -595 64
rect -626 50 -621 55
rect -607 50 -602 55
rect -411 90 -406 95
rect -487 66 -482 71
rect -442 66 -436 71
rect -394 90 -389 95
rect -586 48 -581 53
rect -514 49 -509 54
rect -586 32 -581 37
rect -513 31 -508 36
rect -442 51 -436 56
rect -478 35 -473 40
rect -262 82 -257 88
rect -168 100 -163 105
rect 225 140 230 145
rect 65 111 70 116
rect -319 59 -314 64
rect -337 54 -332 59
rect -359 12 -354 17
rect -273 59 -268 64
rect -299 50 -294 55
rect -280 50 -275 55
rect -84 90 -79 95
rect -160 66 -155 71
rect -115 66 -109 71
rect 15 95 20 100
rect -67 90 -62 95
rect -259 48 -254 53
rect -187 49 -182 54
rect -259 32 -254 37
rect -186 31 -181 36
rect -115 51 -109 56
rect -151 35 -146 40
rect 43 95 48 100
rect 135 106 140 111
rect 206 112 211 117
rect 335 131 340 136
rect 251 111 256 116
rect 322 107 327 112
rect 304 77 309 82
rect 528 226 533 231
rect 697 308 702 313
rect 895 329 901 335
rect 667 242 673 248
rect 573 225 578 230
rect 670 229 675 234
rect 644 221 649 226
rect 692 230 697 235
rect 1012 265 1017 270
rect 989 254 995 260
rect 812 242 818 248
rect 678 185 683 190
rect 816 200 821 205
rect 1172 251 1177 256
rect 1012 222 1017 227
rect 664 174 669 179
rect 359 135 364 140
rect 356 122 361 127
rect 336 105 341 110
rect 450 111 455 116
rect 504 138 509 143
rect 494 120 499 125
rect 337 84 342 89
rect 450 102 455 107
rect 494 107 499 112
rect 450 93 455 98
rect 507 105 512 110
rect 503 93 508 98
rect 975 205 980 210
rect 1082 217 1087 222
rect 1153 223 1158 228
rect 1198 222 1203 227
rect 1269 218 1274 223
rect 585 108 590 113
rect 632 124 637 129
rect 625 110 630 115
rect 594 97 599 102
rect 511 84 516 89
rect 624 98 629 103
rect 639 92 644 97
rect 728 109 733 114
rect 830 127 836 133
rect 829 90 837 98
rect 24 19 29 24
<< labels >>
rlabel metal1 42 854 47 857 4 VDD
rlabel metal1 42 799 47 802 2 GND
rlabel metal1 42 958 46 962 4 VDD
rlabel metal1 42 861 46 865 2 GND
rlabel metal1 146 818 150 822 1 G0
rlabel metal1 335 914 339 918 7 P0
rlabel metal1 351 915 356 918 4 VDD
rlabel metal1 351 860 356 863 2 GND
rlabel metal1 469 915 472 918 4 VDD
rlabel metal1 469 860 472 863 2 GND
rlabel metal1 583 879 587 883 7 C1
rlabel metal1 293 1046 297 1050 4 VDD
rlabel metal1 293 949 297 953 2 GND
rlabel metal1 586 1002 590 1006 7 S0
rlabel metal1 41 674 46 677 4 VDD
rlabel metal1 41 619 46 622 2 GND
rlabel metal1 41 778 45 782 4 VDD
rlabel metal1 41 681 45 685 2 GND
rlabel metal1 145 638 149 642 1 G1
rlabel metal1 334 734 338 738 1 P1
rlabel metal1 357 736 360 739 4 VDD
rlabel metal1 357 681 360 684 2 GND
rlabel metal1 274 829 279 832 4 VDD
rlabel metal1 274 774 279 777 2 GND
rlabel metal1 398 822 401 825 4 VDD
rlabel metal1 426 767 429 770 1 GND
rlabel metal1 531 786 535 790 1 C2
rlabel metal1 173 651 177 655 4 VDD
rlabel metal1 173 554 177 558 2 GND
rlabel metal1 41 420 46 423 4 VDD
rlabel metal1 41 365 46 368 2 GND
rlabel metal1 41 524 45 528 4 VDD
rlabel metal1 41 427 45 431 2 GND
rlabel metal1 362 498 365 501 4 VDD
rlabel metal1 362 443 365 446 2 GND
rlabel metal1 331 480 335 484 1 P2
rlabel metal1 145 384 149 388 1 G2
rlabel metal1 531 499 534 502 4 VDD
rlabel metal1 531 444 534 447 2 GND
rlabel metal1 542 519 545 539 3 VDD
rlabel metal1 531 563 536 566 4 VDD
rlabel metal1 531 508 536 511 2 GND
rlabel metal1 678 511 681 514 4 VDD
rlabel metal1 678 455 681 458 2 GND
rlabel metal1 832 474 836 478 7 C3
rlabel metal1 532 594 536 598 2 GND
rlabel metal1 532 691 536 695 4 VDD
rlabel metal1 42 238 47 241 4 VDD
rlabel metal1 42 183 47 186 2 GND
rlabel metal1 42 342 46 346 4 VDD
rlabel metal1 42 245 46 249 2 GND
rlabel metal1 290 322 293 325 2 GND
rlabel metal1 146 202 150 206 1 G3
rlabel metal1 301 386 306 389 1 VDD
rlabel metal1 426 387 429 390 4 VDD
rlabel metal1 441 332 456 335 1 GND
rlabel metal1 572 387 575 390 4 VDD
rlabel metal1 599 332 604 335 1 GND
rlabel metal1 719 398 722 418 3 VDD
rlabel metal1 708 442 713 445 4 VDD
rlabel metal1 708 387 713 390 2 GND
rlabel metal1 718 366 721 369 4 VDD
rlabel metal1 741 297 749 300 1 GND
rlabel metal1 365 273 369 277 4 VDD
rlabel metal1 365 176 369 180 2 GND
rlabel metal1 335 298 339 302 1 P3
rlabel metal1 43 55 48 58 4 VDD
rlabel metal1 43 0 48 3 2 GND
rlabel metal1 43 159 47 163 4 VDD
rlabel metal1 43 62 47 66 2 GND
rlabel metal1 147 19 151 23 1 G4
rlabel metal1 382 77 386 81 1 VDD
rlabel metal1 470 84 474 88 1 GND
rlabel metal1 290 91 294 95 1 P4
rlabel metal1 508 148 511 151 4 VDD
rlabel metal1 534 84 560 87 1 GND
rlabel metal1 636 84 639 87 2 GND
rlabel metal1 636 139 639 142 4 VDD
rlabel metal1 689 219 692 222 4 VDD
rlabel metal1 712 164 735 167 1 GND
rlabel metal1 846 198 849 218 3 VDD
rlabel metal1 835 242 840 245 4 VDD
rlabel metal1 835 187 840 190 2 GND
rlabel metal1 1034 82 1038 86 1 GND
rlabel metal1 856 81 860 85 1 VDD
rlabel metal1 990 270 994 274 4 VDD
rlabel metal1 990 173 994 177 2 GND
rlabel metal1 890 330 894 334 7 C4
rlabel metal1 -677 981 -674 984 1 VDD
rlabel metal1 -671 867 -667 870 1 GND
rlabel metal1 -692 889 -688 893 3 CLK
rlabel metal1 -677 745 -674 748 1 VDD
rlabel metal1 -671 631 -667 634 1 GND
rlabel metal1 -692 653 -688 657 3 CLK
rlabel metal1 -677 531 -674 534 1 VDD
rlabel metal1 -671 417 -667 420 1 GND
rlabel metal1 -692 439 -688 443 3 CLK
rlabel metal1 -677 292 -674 295 1 VDD
rlabel metal1 -671 178 -667 181 1 GND
rlabel metal1 -692 200 -688 204 3 CLK
rlabel metal1 -677 105 -674 108 1 VDD
rlabel metal1 -671 -9 -667 -6 1 GND
rlabel metal1 -692 13 -688 17 3 CLK
rlabel metal1 -45 976 -40 980 1 B0
rlabel metal1 -45 100 -40 104 1 B4
rlabel metal1 -45 287 -40 291 1 B3
rlabel metal1 -45 526 -40 530 1 B2
rlabel metal1 -45 740 -40 744 1 B1
rlabel metal1 -1336 106 -1333 109 1 VDD
rlabel metal1 -1330 -8 -1326 -5 1 GND
rlabel metal1 -1351 14 -1347 18 3 CLK
rlabel metal1 -1336 293 -1333 296 1 VDD
rlabel metal1 -1330 179 -1326 182 1 GND
rlabel metal1 -1351 201 -1347 205 3 CLK
rlabel metal1 -1336 532 -1333 535 1 VDD
rlabel metal1 -1330 418 -1326 421 1 GND
rlabel metal1 -1351 440 -1347 444 3 CLK
rlabel metal1 -1336 746 -1333 749 1 VDD
rlabel metal1 -1330 632 -1326 635 1 GND
rlabel metal1 -1351 654 -1347 658 3 CLK
rlabel metal1 -1336 985 -1333 988 1 VDD
rlabel metal1 -1330 871 -1326 874 1 GND
rlabel metal1 -1351 893 -1347 897 3 CLK
rlabel metal1 -704 980 -699 984 1 A0
rlabel metal1 -704 741 -699 745 1 A1
rlabel metal1 -704 288 -699 292 1 A3
rlabel metal1 -704 101 -699 105 1 A4
rlabel metal1 -692 944 -688 948 1 B0i
rlabel metal1 -692 708 -688 712 1 B1i
rlabel metal1 -692 494 -688 498 1 B2i
rlabel metal1 -692 255 -688 259 1 B3i
rlabel metal1 -692 68 -688 72 1 B4i
rlabel metal1 -1351 69 -1347 73 3 A4i
rlabel metal1 -1351 256 -1347 260 3 A3i
rlabel metal1 -1351 495 -1347 499 3 A2i
rlabel metal1 -1351 709 -1347 713 3 A1i
rlabel metal1 -1351 948 -1347 952 3 A0i
rlabel metal1 732 727 736 731 1 CLK
rlabel metal1 755 748 758 752 7 GND
rlabel metal1 641 742 644 745 7 VDD
rlabel metal1 874 727 878 731 1 CLK
rlabel metal1 897 748 900 752 7 GND
rlabel metal1 783 742 786 745 7 VDD
rlabel metal1 819 733 823 737 1 S1
rlabel metal1 677 727 681 731 1 S0
rlabel metal1 1014 727 1018 731 1 CLK
rlabel metal1 1037 748 1040 752 7 GND
rlabel metal1 923 742 926 745 7 VDD
rlabel metal1 959 733 963 737 1 S2
rlabel metal1 1159 727 1163 731 1 CLK
rlabel metal1 1182 748 1185 752 7 GND
rlabel metal1 1068 742 1071 745 7 VDD
rlabel metal1 1304 727 1308 731 1 CLK
rlabel metal1 1327 748 1330 752 7 GND
rlabel metal1 1213 742 1216 745 7 VDD
rlabel metal1 1449 727 1453 731 1 CLK
rlabel metal1 1472 748 1475 752 7 GND
rlabel metal1 1358 742 1361 745 7 VDD
rlabel metal1 1104 733 1108 737 1 S3
rlabel metal1 1249 733 1253 737 1 S4
rlabel metal1 1394 733 1398 737 1 Cout
rlabel metal1 645 1374 649 1379 5 S0o
rlabel metal1 787 1374 791 1379 5 S1o
rlabel metal1 927 1374 931 1379 5 S2o
rlabel metal1 1072 1374 1076 1379 5 S3o
rlabel metal1 1217 1374 1221 1379 5 S4o
rlabel metal1 1362 1374 1366 1379 5 Couto
rlabel metal1 -676 1145 -673 1148 1 VDD
rlabel metal1 -670 1031 -666 1034 1 GND
rlabel metal1 -691 1053 -687 1057 3 CLK
rlabel metal1 -44 1140 -39 1144 1 Cin
rlabel metal1 -691 1108 -687 1112 1 Cini
rlabel metal1 -704 527 -699 531 1 A2
<< end >>
