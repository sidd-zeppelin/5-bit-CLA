magic
tech scmos
timestamp 1763746094
<< nwell >>
rect 10 0 102 48
rect 133 21 157 53
<< ntransistor >>
rect 108 35 118 37
rect 108 27 118 29
rect 108 19 118 21
rect 108 11 118 13
rect 144 1 146 11
<< ptransistor >>
rect 16 35 96 37
rect 16 27 96 29
rect 144 27 146 47
rect 16 19 96 21
rect 16 11 96 13
<< ndiffusion >>
rect 108 37 118 38
rect 108 34 118 35
rect 108 29 118 30
rect 108 26 118 27
rect 108 21 118 22
rect 108 18 118 19
rect 108 13 118 14
rect 108 10 118 11
rect 143 1 144 11
rect 146 1 147 11
<< pdiffusion >>
rect 16 37 96 38
rect 16 34 96 35
rect 16 29 96 30
rect 143 27 144 47
rect 146 27 147 47
rect 16 26 96 27
rect 16 21 96 22
rect 16 18 96 19
rect 16 13 96 14
rect 16 10 96 11
<< ndcontact >>
rect 108 38 118 42
rect 108 30 118 34
rect 108 22 118 26
rect 108 14 118 18
rect 108 6 118 10
rect 139 1 143 11
rect 147 1 151 11
<< pdcontact >>
rect 16 38 96 42
rect 16 30 96 34
rect 139 27 143 47
rect 147 27 151 47
rect 16 22 96 26
rect 16 14 96 18
rect 16 6 96 10
<< polysilicon >>
rect 144 47 146 50
rect 7 35 16 37
rect 96 35 108 37
rect 118 35 121 37
rect 7 27 16 29
rect 96 27 108 29
rect 118 27 121 29
rect 7 19 16 21
rect 96 19 108 21
rect 118 19 121 21
rect 7 11 16 13
rect 96 11 108 13
rect 118 11 121 13
rect 144 11 146 27
rect 144 -2 146 1
<< polycontact >>
rect 3 34 7 38
rect 3 26 7 30
rect 3 18 7 22
rect 3 10 7 14
rect 140 14 144 18
<< metal1 >>
rect -1 51 157 54
rect -1 34 3 38
rect -1 26 3 30
rect -1 18 3 22
rect -1 10 3 14
rect 10 10 13 51
rect 101 45 133 48
rect 101 42 104 45
rect 96 38 104 42
rect 118 38 124 42
rect 100 34 104 38
rect 100 30 108 34
rect 100 18 104 30
rect 121 26 124 38
rect 118 22 124 26
rect 100 14 108 18
rect 121 10 124 22
rect 130 18 133 45
rect 139 47 143 51
rect 147 18 151 27
rect 130 14 140 18
rect 147 14 157 18
rect 147 11 151 14
rect 10 6 16 10
rect 118 6 124 10
rect 121 -2 124 6
rect 139 -2 143 1
rect -1 -5 151 -2
<< labels >>
rlabel metal1 -1 10 3 14 3 A
rlabel metal1 -1 18 3 22 3 B
rlabel metal1 -1 26 3 30 3 C
rlabel metal1 -1 34 3 38 3 D
rlabel metal1 153 14 157 18 7 OUT
rlabel metal1 -1 51 2 54 4 VDD
rlabel metal1 -1 -5 2 -2 2 GND
<< end >>
