magic
tech scmos
timestamp 1764589017
<< ntransistor >>
rect 151 34 161 36
rect 151 26 161 28
rect 151 18 161 20
rect 151 10 161 12
rect 151 2 161 4
rect 151 -6 161 -4
<< ptransistor >>
rect 19 34 139 36
rect 19 26 139 28
rect 19 18 139 20
rect 19 10 139 12
rect 19 2 139 4
rect 19 -6 139 -4
<< ndiffusion >>
rect 151 36 161 37
rect 151 33 161 34
rect 151 28 161 29
rect 151 25 161 26
rect 151 20 161 21
rect 151 17 161 18
rect 151 12 161 13
rect 151 9 161 10
rect 151 4 161 5
rect 151 1 161 2
rect 151 -4 161 -3
rect 151 -7 161 -6
<< pdiffusion >>
rect 19 36 139 37
rect 19 33 139 34
rect 19 28 139 29
rect 19 25 139 26
rect 19 20 139 21
rect 19 17 139 18
rect 19 12 139 13
rect 19 9 139 10
rect 19 4 139 5
rect 19 1 139 2
rect 19 -4 139 -3
rect 19 -7 139 -6
<< ndcontact >>
rect 151 37 161 41
rect 151 29 161 33
rect 151 21 161 25
rect 151 13 161 17
rect 151 5 161 9
rect 151 -3 161 1
rect 151 -11 161 -7
<< pdcontact >>
rect 19 37 139 41
rect 19 29 139 33
rect 19 21 139 25
rect 19 13 139 17
rect 19 5 139 9
rect 19 -3 139 1
rect 19 -11 139 -7
<< polysilicon >>
rect 8 34 19 36
rect 139 34 151 36
rect 161 34 164 36
rect 8 26 19 28
rect 139 26 151 28
rect 161 26 164 28
rect 8 18 19 20
rect 139 18 151 20
rect 161 18 164 20
rect 8 10 19 12
rect 139 10 151 12
rect 161 10 164 12
rect 8 2 19 4
rect 139 2 151 4
rect 161 2 164 4
rect 8 -6 19 -4
rect 139 -6 151 -4
rect 161 -6 164 -4
<< polycontact >>
rect 4 33 8 37
rect 4 25 8 29
rect 4 17 8 21
rect 4 9 8 13
rect 4 1 8 5
rect 4 -7 8 -3
<< metal1 >>
rect 142 45 172 49
rect 142 41 146 45
rect 0 33 4 37
rect 0 25 4 29
rect 0 17 4 21
rect 0 9 4 13
rect 0 1 4 5
rect 0 -7 4 -3
rect 11 -7 15 41
rect 139 37 146 41
rect 161 37 168 41
rect 142 33 146 37
rect 142 29 151 33
rect 142 17 146 29
rect 164 25 168 37
rect 161 21 168 25
rect 142 13 151 17
rect 142 1 146 13
rect 164 9 168 21
rect 161 5 168 9
rect 142 -3 151 1
rect 164 -7 168 5
rect 11 -11 19 -7
rect 161 -11 168 -7
<< labels >>
rlabel metal1 11 -11 15 41 3 VDD
rlabel metal1 164 -11 168 41 7 GND
rlabel metal1 168 45 172 49 6 OUT
rlabel metal1 0 -7 4 -3 3 A
rlabel metal1 0 1 4 5 3 B
rlabel metal1 0 9 4 13 3 C
rlabel metal1 0 17 4 21 3 D
rlabel metal1 0 25 4 29 3 E
rlabel metal1 0 33 4 37 3 F
<< end >>
