magic
tech scmos
timestamp 1763748553
<< nwell >>
rect 11 0 123 56
rect 152 33 176 65
<< ntransistor >>
rect 129 43 139 45
rect 129 35 139 37
rect 129 27 139 29
rect 129 19 139 21
rect 163 13 165 23
rect 129 11 139 13
<< ptransistor >>
rect 17 43 117 45
rect 163 39 165 59
rect 17 35 117 37
rect 17 27 117 29
rect 17 19 117 21
rect 17 11 117 13
<< ndiffusion >>
rect 129 45 139 46
rect 129 42 139 43
rect 129 37 139 38
rect 129 34 139 35
rect 129 29 139 30
rect 129 26 139 27
rect 129 21 139 22
rect 129 18 139 19
rect 129 13 139 14
rect 162 13 163 23
rect 165 13 166 23
rect 129 10 139 11
<< pdiffusion >>
rect 17 45 117 46
rect 17 42 117 43
rect 17 37 117 38
rect 162 39 163 59
rect 165 39 166 59
rect 17 34 117 35
rect 17 29 117 30
rect 17 26 117 27
rect 17 21 117 22
rect 17 18 117 19
rect 17 13 117 14
rect 17 10 117 11
<< ndcontact >>
rect 129 46 139 50
rect 129 38 139 42
rect 129 30 139 34
rect 129 22 139 26
rect 129 14 139 18
rect 158 13 162 23
rect 166 13 170 23
rect 129 6 139 10
<< pdcontact >>
rect 17 46 117 50
rect 17 38 117 42
rect 158 39 162 59
rect 166 39 170 59
rect 17 30 117 34
rect 17 22 117 26
rect 17 14 117 18
rect 17 6 117 10
<< polysilicon >>
rect 163 59 165 62
rect 8 43 17 45
rect 117 43 129 45
rect 139 43 142 45
rect 8 35 17 37
rect 117 35 129 37
rect 139 35 142 37
rect 8 27 17 29
rect 117 27 129 29
rect 139 27 142 29
rect 163 23 165 39
rect 8 19 17 21
rect 117 19 129 21
rect 139 19 142 21
rect 8 11 17 13
rect 117 11 129 13
rect 139 11 142 13
rect 163 10 165 13
<< polycontact >>
rect 4 42 8 46
rect 4 34 8 38
rect 4 26 8 30
rect 4 18 8 22
rect 159 26 163 30
rect 4 10 8 14
<< metal1 >>
rect 0 62 176 65
rect 0 42 4 46
rect 0 34 4 38
rect 0 26 4 30
rect 0 18 4 22
rect 0 10 4 14
rect 11 10 14 62
rect 158 59 162 62
rect 123 53 152 56
rect 123 50 126 53
rect 117 46 129 50
rect 122 34 126 46
rect 142 42 145 50
rect 139 38 145 42
rect 122 30 129 34
rect 122 18 126 30
rect 142 26 145 38
rect 149 30 152 53
rect 166 30 170 39
rect 149 26 159 30
rect 166 26 176 30
rect 139 22 145 26
rect 166 23 170 26
rect 122 14 129 18
rect 142 10 145 22
rect 11 6 17 10
rect 139 9 145 10
rect 158 9 162 13
rect 139 6 162 9
rect 11 0 14 6
rect 142 -4 145 6
rect 0 -7 145 -4
<< labels >>
rlabel metal1 0 10 4 14 3 A
rlabel metal1 0 18 4 22 3 B
rlabel metal1 0 26 4 30 3 C
rlabel metal1 0 34 4 38 3 D
rlabel metal1 0 42 4 46 3 E
rlabel metal1 172 26 176 30 7 OUT
rlabel metal1 0 -7 3 -4 2 GND
rlabel metal1 0 62 3 65 4 VDD
<< end >>
