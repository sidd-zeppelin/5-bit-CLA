* SPICE3 file created from NAND5.ext - technology: scmos

.option scale=0.09u

M1000 OUT C VDD w_n6_31# cmosp w=20 l=2
+  ad=340 pd=154 as=340 ps=154
M1001 a_31_0# D a_23_0# Gnd cmosn w=25 l=2
+  ad=150 pd=62 as=150 ps=62
M1002 VDD D OUT w_n6_31# cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1003 a_15_0# B a_7_0# Gnd cmosn w=25 l=2
+  ad=150 pd=62 as=150 ps=62
M1004 OUT A VDD w_n6_31# cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1005 VDD B OUT w_n6_31# cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
M1006 a_7_0# A GND Gnd cmosn w=25 l=2
+  ad=0 pd=0 as=125 ps=60
M1007 OUT E a_31_0# Gnd cmosn w=25 l=2
+  ad=125 pd=60 as=0 ps=0
M1008 a_23_0# C a_15_0# Gnd cmosn w=25 l=2
+  ad=0 pd=0 as=0 ps=0
M1009 OUT E VDD w_n6_31# cmosp w=20 l=2
+  ad=0 pd=0 as=0 ps=0
