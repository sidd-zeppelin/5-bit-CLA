magic
tech scmos
timestamp 1764588226
<< nwell >>
rect 11 0 34 64
rect 93 33 117 65
<< ntransistor >>
rect 42 51 72 53
rect 42 43 72 45
rect 42 35 72 37
rect 42 27 72 29
rect 42 19 72 21
rect 104 13 106 23
rect 42 11 72 13
<< ptransistor >>
rect 18 51 28 53
rect 18 43 28 45
rect 104 39 106 59
rect 18 35 28 37
rect 18 27 28 29
rect 18 19 28 21
rect 18 11 28 13
<< ndiffusion >>
rect 42 53 72 54
rect 42 50 72 51
rect 42 45 72 46
rect 42 42 72 43
rect 42 37 72 38
rect 42 34 72 35
rect 42 29 72 30
rect 42 26 72 27
rect 42 21 72 22
rect 42 18 72 19
rect 42 13 72 14
rect 103 13 104 23
rect 106 13 107 23
rect 42 10 72 11
<< pdiffusion >>
rect 18 53 28 54
rect 18 50 28 51
rect 18 45 28 46
rect 18 42 28 43
rect 18 37 28 38
rect 103 39 104 59
rect 106 39 107 59
rect 18 34 28 35
rect 18 29 28 30
rect 18 26 28 27
rect 18 21 28 22
rect 18 18 28 19
rect 18 13 28 14
rect 18 10 28 11
<< ndcontact >>
rect 42 54 72 58
rect 42 46 72 50
rect 42 38 72 42
rect 42 30 72 34
rect 42 22 72 26
rect 42 14 72 18
rect 99 13 103 23
rect 107 13 111 23
rect 42 6 72 10
<< pdcontact >>
rect 18 54 28 58
rect 18 46 28 50
rect 18 38 28 42
rect 99 39 103 59
rect 107 39 111 59
rect 18 30 28 34
rect 18 22 28 26
rect 18 14 28 18
rect 18 6 28 10
<< polysilicon >>
rect 104 59 106 62
rect 8 51 18 53
rect 28 51 42 53
rect 72 51 75 53
rect 8 43 18 45
rect 28 43 42 45
rect 72 43 75 45
rect 8 35 18 37
rect 28 35 42 37
rect 72 35 75 37
rect 8 27 18 29
rect 28 27 42 29
rect 72 27 75 29
rect 104 23 106 39
rect 8 19 18 21
rect 28 19 42 21
rect 72 19 75 21
rect 8 11 18 13
rect 28 11 42 13
rect 72 11 75 13
rect 104 10 106 13
<< polycontact >>
rect 4 50 8 54
rect 4 42 8 46
rect 4 34 8 38
rect 4 26 8 30
rect 4 18 8 22
rect 100 26 104 30
rect 4 10 8 14
<< metal1 >>
rect 11 73 97 77
rect 11 58 15 73
rect 93 65 97 73
rect 34 61 90 65
rect 93 62 103 65
rect 34 58 38 61
rect 11 54 18 58
rect 34 54 42 58
rect 0 50 4 54
rect 0 42 4 46
rect 11 42 15 54
rect 34 50 38 54
rect 28 46 38 50
rect 11 38 18 42
rect 0 34 4 38
rect 0 26 4 30
rect 11 26 15 38
rect 34 34 38 46
rect 28 30 38 34
rect 86 30 90 61
rect 99 59 103 62
rect 107 30 111 39
rect 11 22 18 26
rect 0 18 4 22
rect 0 10 4 14
rect 11 10 15 22
rect 34 18 38 30
rect 86 26 100 30
rect 107 26 117 30
rect 107 23 111 26
rect 28 14 38 18
rect 99 10 103 13
rect 11 6 18 10
rect 72 7 103 10
rect 72 6 75 7
rect 11 0 15 6
<< labels >>
rlabel metal1 0 10 4 14 3 A
rlabel metal1 0 18 4 22 3 B
rlabel metal1 0 26 4 30 3 C
rlabel metal1 0 34 4 38 3 D
rlabel metal1 0 42 4 46 3 E
rlabel metal1 0 50 4 54 3 F
rlabel metal1 113 26 117 30 7 OUT
rlabel metal1 11 0 15 4 1 VDD
rlabel metal1 99 7 103 11 1 GND
<< end >>
