* SPICE3 file created from OR4.ext - technology: scmos

.option scale=0.09u

M1000 GND D a_16_37# Gnd cmosn w=10 l=2
+  ad=210 pd=122 as=120 ps=64
M1001 OUT a_16_37# GND Gnd cmosn w=10 l=2
+  ad=50 pd=30 as=0 ps=0
M1002 a_16_21# B a_16_13# w_10_0# cmosp w=80 l=2
+  ad=480 pd=172 as=480 ps=172
M1003 GND B a_16_37# Gnd cmosn w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1004 a_16_29# C a_16_21# w_10_0# cmosp w=80 l=2
+  ad=480 pd=172 as=0 ps=0
M1005 a_16_13# A VDD w_10_0# cmosp w=80 l=2
+  ad=0 pd=0 as=500 ps=220
M1006 OUT a_16_37# VDD w_133_21# cmosp w=20 l=2
+  ad=100 pd=50 as=0 ps=0
M1007 a_16_37# C GND Gnd cmosn w=10 l=2
+  ad=0 pd=0 as=0 ps=0
M1008 a_16_37# D a_16_29# w_10_0# cmosp w=80 l=2
+  ad=400 pd=170 as=0 ps=0
M1009 a_16_37# A GND Gnd cmosn w=10 l=2
+  ad=0 pd=0 as=0 ps=0
C0 w_10_0# Gnd 4.44fF
