* NGSPICE file created from cla.ext - technology: scmos

.global Vdd Gnd 


* Top level circuit cla

M1000 a_693_n302# G2 GND Gnd cmosn w=0.9u l=0.18u
+  ad=0.972p pd=5.76u as=51.9615p ps=296.82u
M1001 a_486_n609# C3 VDD w_480_n622# cmosp w=1.8u l=0.18u
+  ad=0.972p pd=4.68u as=104.004p ps=563.76u
M1002 a_163_132# a_72_98# VDD w_157_119# cmosp w=1.8u l=0.18u
+  ad=0.972p pd=4.68u as=0p ps=0u
M1003 a_400_n7# a_372_n97# GND Gnd cmosn w=0.9u l=0.18u
+  ad=0.405p pd=2.7u as=0p ps=0u
M1004 a_294_n175# a_203_n209# VDD w_288_n188# cmosp w=1.8u l=0.18u
+  ad=0.972p pd=4.68u as=0p ps=0u
M1005 VDD P3 a_395_n587# w_389_n600# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1006 G2 a_56_n416# GND Gnd cmosn w=0.9u l=0.18u
+  ad=0.405p pd=2.7u as=0p ps=0u
M1007 GND a_562_n169# a_689_n191# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1008 GND a_203_n209# a_330_n231# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1009 a_163_n484# a_72_n518# VDD w_157_n497# cmosp w=1.8u l=0.18u
+  ad=0.972p pd=4.68u as=0p ps=0u
M1010 a_390_n462# a_305_n461# GND Gnd cmosn w=0.9u l=0.18u
+  ad=0.405p pd=2.7u as=0p ps=0u
M1011 a_162_n358# B2 VDD w_156_n371# cmosp w=1.8u l=0.18u
+  ad=0.972p pd=4.68u as=0p ps=0u
M1012 a_473_n435# P1 a_473_n443# Gnd cmosn w=3.6u l=0.18u
+  ad=1.944p pd=8.28u as=1.944p ps=8.28u
M1013 a_441_n451# P1 VDD w_435_n464# cmosp w=1.8u l=0.18u
+  ad=1.944p pd=9.36u as=0p ps=0u
M1014 a_89_n416# B2 GND Gnd cmosn w=1.8u l=0.18u
+  ad=0.972p pd=4.68u as=0p ps=0u
M1015 VDD A2 a_56_n416# w_50_n429# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1016 a_587_n446# G1 a_619_n438# Gnd cmosn w=2.7u l=0.18u
+  ad=1.215p pd=6.3u as=1.458p ps=6.48u
M1017 VDD A2 a_162_n302# w_156_n315# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1018 GND Cin a_450_220# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1019 a_635_n349# a_546_n334# VDD w_622_n329# cmosp w=1.8u l=0.18u
+  ad=0.81p pd=4.5u as=0p ps=0u
M1020 GND a_486_n553# a_618_n587# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1021 a_400_n7# a_372_n97# VDD w_448_n92# cmosp w=1.8u l=0.18u
+  ad=0.81p pd=4.5u as=0p ps=0u
M1022 S2 a_653_n191# VDD w_743_n182# cmosp w=1.8u l=0.18u
+  ad=0.972p pd=4.68u as=0p ps=0u
M1023 a_693_n326# G2 VDD w_687_n339# cmosp w=7.2u l=0.18u
+  ad=3.888p pd=15.48u as=0p ps=0u
M1024 a_450_164# P0 a_414_164# Gnd cmosn w=1.8u l=0.18u
+  ad=0.972p pd=4.68u as=0.81p ps=4.5u
M1025 a_369_n19# a_289_n7# GND Gnd cmosn w=0.9u l=0.18u
+  ad=0.405p pd=2.7u as=0p ps=0u
M1026 a_372_n97# P1 a_404_n89# Gnd cmosn w=2.7u l=0.18u
+  ad=1.215p pd=6.3u as=1.458p ps=6.48u
M1027 VDD a_203_n209# a_294_n231# w_288_n244# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1028 a_693_n302# a_476_n350# GND Gnd cmosn w=0.9u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1029 GND Cin a_359_186# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1030 P0 a_163_76# VDD w_253_85# cmosp w=1.8u l=0.18u
+  ad=0.972p pd=4.68u as=0p ps=0u
M1031 GND P3 a_522_n553# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1032 VDD a_72_n518# a_163_n540# w_157_n553# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1033 G2 a_56_n416# VDD w_123_n408# cmosp w=1.8u l=0.18u
+  ad=0.81p pd=4.5u as=0p ps=0u
M1034 a_653_n135# a_562_n169# VDD w_647_n148# cmosp w=1.8u l=0.18u
+  ad=0.972p pd=4.68u as=0p ps=0u
M1035 a_203_n209# C1 VDD w_197_n222# cmosp w=1.8u l=0.18u
+  ad=0.972p pd=4.68u as=0p ps=0u
M1036 a_484_86# G0 GND Gnd cmosn w=0.9u l=0.18u
+  ad=0.486p pd=2.88u as=0p ps=0u
M1037 VDD a_162_n48# P1 w_252_n95# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1038 a_56_n162# B1 VDD w_50_n175# cmosp w=1.8u l=0.18u
+  ad=0.972p pd=4.68u as=0p ps=0u
M1039 a_413_4# a_369_n19# a_413_n4# w_407_n25# cmosp w=5.4u l=0.18u
+  ad=2.43p pd=11.7u as=2.916p ps=11.88u
M1040 G1 a_56_n162# VDD w_123_n154# cmosp w=1.8u l=0.18u
+  ad=0.81p pd=4.5u as=0p ps=0u
M1041 a_723_n394# P3 VDD w_717_n407# cmosp w=1.8u l=0.18u
+  ad=0.972p pd=4.68u as=0p ps=0u
M1042 a_294_n336# a_162_n358# P2 Gnd cmosn w=1.8u l=0.18u
+  ad=0.972p pd=4.68u as=0.81p ps=4.5u
M1043 a_108_n518# B3 a_72_n518# Gnd cmosn w=1.8u l=0.18u
+  ad=0.972p pd=4.68u as=0.81p ps=4.5u
M1044 a_546_n334# G0 a_578_n326# Gnd cmosn w=2.7u l=0.18u
+  ad=1.215p pd=6.3u as=1.458p ps=6.48u
M1045 a_733_n450# G3 GND Gnd cmosn w=0.9u l=0.18u
+  ad=1.377p pd=8.46u as=0p ps=0u
M1046 a_733_n466# a_540_n461# a_733_n474# w_727_n495# cmosp w=9u l=0.18u
+  ad=4.86p pd=19.08u as=4.86p ps=19.08u
M1047 a_57_18# B0 VDD w_51_5# cmosp w=1.8u l=0.18u
+  ad=0.972p pd=4.68u as=0p ps=0u
M1048 a_546_n334# G0 VDD w_540_n347# cmosp w=1.8u l=0.18u
+  ad=1.782p pd=9.18u as=0p ps=0u
M1049 VDD a_562_n169# a_653_n191# w_647_n204# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1050 VDD a_163_132# P0 w_253_85# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1051 a_198_n48# a_71_n82# a_162_n48# Gnd cmosn w=1.8u l=0.18u
+  ad=0.972p pd=4.68u as=0.81p ps=4.5u
M1052 a_409_n340# P2 GND Gnd cmosn w=3.6u l=0.18u
+  ad=1.944p pd=8.28u as=0p ps=0u
M1053 a_337_n461# P3 GND Gnd cmosn w=2.25u l=0.18u
+  ad=1.215p pd=5.58u as=0p ps=0u
M1054 a_720_n453# a_723_n394# GND Gnd cmosn w=0.9u l=0.18u
+  ad=0.405p pd=2.7u as=0p ps=0u
M1055 a_198_n302# a_71_n336# a_162_n302# Gnd cmosn w=1.8u l=0.18u
+  ad=0.972p pd=4.68u as=0.81p ps=4.5u
M1056 C3 a_693_n302# GND Gnd cmosn w=0.9u l=0.18u
+  ad=0.405p pd=2.7u as=0p ps=0u
M1057 a_305_n461# P3 VDD w_299_n474# cmosp w=1.8u l=0.18u
+  ad=2.754p pd=13.86u as=0p ps=0u
M1058 C2 a_413_4# GND Gnd cmosn w=0.9u l=0.18u
+  ad=0.405p pd=2.7u as=0p ps=0u
M1059 a_199_n540# B3 a_163_n540# Gnd cmosn w=1.8u l=0.18u
+  ad=0.972p pd=4.68u as=0.81p ps=4.5u
M1060 VDD P3 a_486_n553# w_480_n566# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1061 VDD Cin a_323_186# w_317_173# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1062 GND A2 a_107_n336# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1063 a_693_n310# a_476_n350# a_693_n318# w_687_n339# cmosp w=7.2u l=0.18u
+  ad=3.888p pd=15.48u as=3.888p ps=15.48u
M1064 a_90_18# B0 GND Gnd cmosn w=1.8u l=0.18u
+  ad=0.972p pd=4.68u as=0p ps=0u
M1065 C4 a_733_n450# VDD w_868_n462# cmosp w=1.8u l=0.18u
+  ad=0.81p pd=4.5u as=0p ps=0u
M1066 GND a_72_98# a_199_76# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1067 P3 a_163_n540# VDD w_253_n531# cmosp w=1.8u l=0.18u
+  ad=0.972p pd=4.68u as=0p ps=0u
M1068 GND a_163_n484# a_295_n518# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1069 a_377_n340# P0 VDD w_371_n353# cmosp w=1.8u l=0.18u
+  ad=1.944p pd=9.36u as=0p ps=0u
M1070 VDD a_323_186# a_414_164# w_408_151# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1071 GND a_676_n461# a_733_n450# Gnd cmosn w=0.9u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1072 VDD P2 a_587_n446# w_581_n459# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=1.782p ps=9.18u
M1073 GND a_71_n82# a_198_n104# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1074 GND a_162_n48# a_294_n82# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1075 GND a_71_n336# a_198_n358# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1076 a_372_n97# Cin VDD w_366_n110# cmosp w=1.8u l=0.18u
+  ad=1.782p pd=9.18u as=0p ps=0u
M1077 a_626_n285# a_546_n273# VDD w_613_n265# cmosp w=1.8u l=0.18u
+  ad=0.81p pd=4.5u as=0p ps=0u
M1078 a_377_n340# Cin a_409_n324# Gnd cmosn w=3.6u l=0.18u
+  ad=1.62p pd=8.1u as=1.944p ps=8.28u
M1079 a_337_n437# P0 a_337_n445# Gnd cmosn w=2.25u l=0.18u
+  ad=1.215p pd=5.58u as=1.215p ps=5.58u
M1080 G0 a_57_18# VDD w_124_26# cmosp w=1.8u l=0.18u
+  ad=0.81p pd=4.5u as=0p ps=0u
M1081 G0 a_57_18# GND Gnd cmosn w=0.9u l=0.18u
+  ad=0.405p pd=2.7u as=0p ps=0u
M1082 a_689_n191# P2 a_653_n191# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.81p ps=4.5u
M1083 a_330_n231# C1 a_294_n231# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.81p ps=4.5u
M1084 a_546_n273# G1 a_579_n273# Gnd cmosn w=1.8u l=0.18u
+  ad=0.81p pd=4.5u as=0.972p ps=4.68u
M1085 VDD P0 a_305_n461# w_299_n474# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1086 a_413_4# G1 GND Gnd cmosn w=0.9u l=0.18u
+  ad=0.891p pd=5.58u as=0p ps=0u
M1087 VDD G0 a_289_n7# w_283_n20# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1088 a_162_n48# a_71_n82# VDD w_156_n61# cmosp w=1.8u l=0.18u
+  ad=0.972p pd=4.68u as=0p ps=0u
M1089 VDD a_162_n302# P2 w_252_n349# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1090 a_72_98# B0 VDD w_66_85# cmosp w=1.8u l=0.18u
+  ad=0.972p pd=4.68u as=0p ps=0u
M1091 a_163_76# B0 VDD w_157_63# cmosp w=1.8u l=0.18u
+  ad=0.972p pd=4.68u as=0p ps=0u
M1092 GND a_653_n135# a_785_n169# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1093 a_733_n450# a_720_n453# a_733_n458# w_727_n495# cmosp w=9u l=0.18u
+  ad=4.05p pd=18.9u as=4.86p ps=19.08u
M1094 a_366_79# P0 VDD w_360_66# cmosp w=1.8u l=0.18u
+  ad=0.972p pd=4.68u as=0p ps=0u
M1095 a_540_n461# a_441_n451# GND Gnd cmosn w=0.9u l=0.18u
+  ad=0.405p pd=2.7u as=0p ps=0u
M1096 a_473_n443# P2 a_473_n451# Gnd cmosn w=3.6u l=0.18u
+  ad=0p pd=0u as=1.944p ps=8.28u
M1097 VDD P2 a_441_n451# w_435_n464# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1098 a_56_n416# B2 VDD w_50_n429# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1099 GND a_163_132# a_295_98# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1100 C3 a_693_n302# VDD w_810_n318# cmosp w=1.8u l=0.18u
+  ad=0.81p pd=4.5u as=0p ps=0u
M1101 GND a_400_n7# a_413_4# Gnd cmosn w=0.9u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1102 GND C2 a_598_n169# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1103 a_90_n598# B3 GND Gnd cmosn w=1.8u l=0.18u
+  ad=0.972p pd=4.68u as=0p ps=0u
M1104 a_390_n462# a_305_n461# VDD w_377_n442# cmosp w=1.8u l=0.18u
+  ad=0.81p pd=4.5u as=0p ps=0u
M1105 C1 a_484_86# VDD w_561_87# cmosp w=1.8u l=0.18u
+  ad=0.81p pd=4.5u as=0p ps=0u
M1106 VDD a_71_n82# a_162_n104# w_156_n117# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1107 VDD A3 a_57_n598# w_51_n611# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1108 a_546_186# a_414_164# S0 Gnd cmosn w=1.8u l=0.18u
+  ad=0.972p pd=4.68u as=0.81p ps=4.5u
M1109 C1 a_484_86# GND Gnd cmosn w=0.9u l=0.18u
+  ad=0.405p pd=2.7u as=0p ps=0u
M1110 GND a_323_186# a_450_164# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1111 a_404_n89# P0 a_404_n97# Gnd cmosn w=2.7u l=0.18u
+  ad=0p pd=0u as=1.458p ps=6.48u
M1112 a_294_n231# C1 VDD w_288_n244# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1113 a_72_n518# B3 VDD w_66_n531# cmosp w=1.8u l=0.18u
+  ad=0.972p pd=4.68u as=0p ps=0u
M1114 a_162_n302# a_71_n336# VDD w_156_n315# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1115 a_431_n587# C3 a_395_n587# Gnd cmosn w=1.8u l=0.18u
+  ad=0.972p pd=4.68u as=0.81p ps=4.5u
M1116 GND A0 a_199_132# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1117 a_522_n553# a_395_n587# a_486_n553# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.81p ps=4.5u
M1118 a_163_n540# B3 VDD w_157_n553# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1119 a_399_79# P0 GND Gnd cmosn w=1.8u l=0.18u
+  ad=0.972p pd=4.68u as=0p ps=0u
M1120 GND a_446_67# a_484_86# Gnd cmosn w=0.9u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1121 a_289_n7# P1 VDD w_283_n20# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1122 P1 a_162_n104# VDD w_252_n95# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1123 VDD a_294_n175# S1 w_384_n222# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1124 a_372_n97# P1 VDD w_366_n110# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1125 GND A1 a_107_n82# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1126 VDD A2 a_71_n336# w_65_n349# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1127 a_676_n461# a_587_n446# GND Gnd cmosn w=0.9u l=0.18u
+  ad=0.405p pd=2.7u as=0p ps=0u
M1128 a_484_78# G0 VDD w_478_65# cmosp w=3.6u l=0.18u
+  ad=1.944p pd=8.28u as=0p ps=0u
M1129 VDD A1 a_71_n82# w_65_n95# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1130 a_413_n4# a_400_n7# a_413_n12# w_407_n25# cmosp w=5.4u l=0.18u
+  ad=0p pd=0u as=2.916p ps=11.88u
M1131 a_578_n326# P1 a_578_n334# Gnd cmosn w=2.7u l=0.18u
+  ad=0p pd=0u as=1.458p ps=6.48u
M1132 S3 a_486_n609# VDD w_576_n600# cmosp w=1.8u l=0.18u
+  ad=0.972p pd=4.68u as=0p ps=0u
M1133 a_733_n474# a_390_n462# a_733_n482# w_727_n495# cmosp w=9u l=0.18u
+  ad=0p pd=0u as=4.86p ps=19.08u
M1134 GND A3 a_199_n484# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1135 VDD a_71_n336# a_162_n358# w_156_n371# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1136 VDD A0 a_57_18# w_51_5# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1137 VDD P1 a_546_n334# w_540_n347# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1138 a_653_n191# P2 VDD w_647_n204# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1139 S0 a_414_164# VDD w_504_173# cmosp w=1.8u l=0.18u
+  ad=0.972p pd=4.68u as=0p ps=0u
M1140 GND A0 a_108_98# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1141 a_56_n162# A1 a_89_n162# Gnd cmosn w=1.8u l=0.18u
+  ad=0.81p pd=4.5u as=0.972p ps=4.68u
M1142 VDD A0 a_163_132# w_157_119# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1143 a_395_n587# C3 VDD w_389_n600# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1144 a_486_n553# a_395_n587# VDD w_480_n566# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1145 a_720_n453# a_723_n394# VDD w_790_n386# cmosp w=1.8u l=0.18u
+  ad=0.81p pd=4.5u as=0p ps=0u
M1146 a_107_n336# B2 a_71_n336# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.81p ps=4.5u
M1147 a_476_n350# a_377_n340# GND Gnd cmosn w=0.9u l=0.18u
+  ad=0.405p pd=2.7u as=0p ps=0u
M1148 GND a_395_n587# a_522_n609# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1149 a_723_n394# G2 a_756_n394# Gnd cmosn w=1.8u l=0.18u
+  ad=0.81p pd=4.5u as=0.972p ps=4.68u
M1150 VDD A0 a_72_98# w_66_85# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1151 a_57_18# A0 a_90_18# Gnd cmosn w=1.8u l=0.18u
+  ad=0.81p pd=4.5u as=0p ps=0u
M1152 a_289_n7# G0 a_322_n7# Gnd cmosn w=1.8u l=0.18u
+  ad=0.81p pd=4.5u as=0.972p ps=4.68u
M1153 GND P1 a_330_n175# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1154 VDD P1 a_377_n340# w_371_n353# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1155 VDD C2 a_562_n169# w_556_n182# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1156 a_733_n450# a_540_n461# GND Gnd cmosn w=0.9u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1157 a_587_n446# P3 VDD w_581_n459# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1158 GND a_294_n175# a_426_n209# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1159 a_294_n82# a_162_n104# P1 Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.81p ps=4.5u
M1160 a_413_n12# G1 VDD w_407_n25# cmosp w=5.4u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1161 a_409_n324# P0 a_409_n332# Gnd cmosn w=3.6u l=0.18u
+  ad=0p pd=0u as=1.944p ps=8.28u
M1162 a_619_n438# P2 a_619_n446# Gnd cmosn w=2.7u l=0.18u
+  ad=0p pd=0u as=1.458p ps=6.48u
M1163 a_337_n445# P1 a_337_n453# Gnd cmosn w=2.25u l=0.18u
+  ad=0p pd=0u as=1.215p ps=5.58u
M1164 VDD G1 a_546_n273# w_540_n286# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1165 a_579_n273# P2 GND Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1166 a_305_n461# P1 VDD w_299_n474# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1167 GND C2 a_689_n135# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1168 GND P1 a_239_n209# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.972p ps=4.68u
M1169 P2 a_162_n358# VDD w_252_n349# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1170 G3 a_57_n598# GND Gnd cmosn w=0.9u l=0.18u
+  ad=0.405p pd=2.7u as=0p ps=0u
M1171 a_414_220# a_323_186# VDD w_408_207# cmosp w=1.8u l=0.18u
+  ad=0.972p pd=4.68u as=0p ps=0u
M1172 VDD a_72_98# a_163_76# w_157_63# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1173 a_369_n19# a_289_n7# VDD w_356_1# cmosp w=1.8u l=0.18u
+  ad=0.81p pd=4.5u as=0p ps=0u
M1174 a_618_n587# a_486_n609# S3 Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.81p ps=4.5u
M1175 GND A3 a_108_n518# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1176 a_785_n169# a_653_n191# S2 Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.81p ps=4.5u
M1177 VDD Cin a_366_79# w_360_66# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1178 a_413_4# a_369_n19# GND Gnd cmosn w=0.9u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1179 a_473_n451# P3 GND Gnd cmosn w=3.6u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1180 a_441_n451# P3 VDD w_435_n464# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1181 GND A1 a_198_n48# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1182 GND a_635_n349# a_693_n302# Gnd cmosn w=0.9u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1183 VDD a_395_n587# a_486_n609# w_480_n622# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1184 a_198_n104# B1 a_162_n104# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.81p ps=4.5u
M1185 a_598_n169# P2 a_562_n169# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.81p ps=4.5u
M1186 VDD P1 a_294_n175# w_288_n188# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1187 a_476_n350# a_377_n340# VDD w_463_n330# cmosp w=1.8u l=0.18u
+  ad=0.81p pd=4.5u as=0p ps=0u
M1188 VDD A3 a_163_n484# w_157_n497# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1189 GND a_414_220# a_546_186# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1190 a_295_98# a_163_76# P0 Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.81p ps=4.5u
M1191 G3 a_57_n598# VDD w_124_n590# cmosp w=1.8u l=0.18u
+  ad=0.81p pd=4.5u as=0p ps=0u
M1192 VDD a_163_n484# P3 w_253_n531# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1193 a_540_n461# a_441_n451# VDD w_527_n441# cmosp w=1.8u l=0.18u
+  ad=0.81p pd=4.5u as=0p ps=0u
M1194 a_733_n450# a_720_n453# GND Gnd cmosn w=0.9u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1195 a_587_n446# G1 VDD w_581_n459# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1196 a_441_n451# G0 a_473_n435# Gnd cmosn w=3.6u l=0.18u
+  ad=1.62p pd=8.1u as=0p ps=0u
M1197 a_366_79# Cin a_399_79# Gnd cmosn w=1.8u l=0.18u
+  ad=0.81p pd=4.5u as=0p ps=0u
M1198 VDD G0 a_441_n451# w_435_n464# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1199 a_56_n416# A2 a_89_n416# Gnd cmosn w=1.8u l=0.18u
+  ad=0.81p pd=4.5u as=0p ps=0u
M1200 S1 a_294_n231# VDD w_384_n222# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1201 a_305_n461# Cin a_337_n437# Gnd cmosn w=2.25u l=0.18u
+  ad=1.0125p pd=5.4u as=0p ps=0u
M1202 a_322_n7# P1 GND Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1203 VDD P0 a_372_n97# w_366_n110# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1204 a_305_n461# Cin VDD w_299_n474# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1205 a_107_n82# B1 a_71_n82# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.81p ps=4.5u
M1206 VDD A1 a_162_n48# w_156_n61# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1207 a_450_220# a_323_186# a_414_220# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.81p ps=4.5u
M1208 G1 a_56_n162# GND Gnd cmosn w=0.9u l=0.18u
+  ad=0.405p pd=2.7u as=0p ps=0u
M1209 a_71_n336# B2 VDD w_65_n349# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1210 a_484_86# a_446_67# a_484_78# w_478_65# cmosp w=3.6u l=0.18u
+  ad=1.62p pd=8.1u as=0p ps=0u
M1211 a_71_n82# B1 VDD w_65_n95# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1212 VDD a_653_n135# S2 w_743_n182# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1213 a_693_n318# a_635_n349# a_693_n326# w_687_n339# cmosp w=7.2u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1214 a_578_n334# P2 GND Gnd cmosn w=2.7u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1215 a_733_n482# G3 VDD w_727_n495# cmosp w=9u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1216 a_199_n484# a_72_n518# a_163_n484# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.81p ps=4.5u
M1217 C2 a_413_4# VDD w_509_n6# cmosp w=1.8u l=0.18u
+  ad=0.81p pd=4.5u as=0p ps=0u
M1218 a_546_n334# P2 VDD w_540_n347# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1219 a_295_n518# a_163_n540# P3 Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.81p ps=4.5u
M1220 a_446_67# a_366_79# VDD w_433_87# cmosp w=1.8u l=0.18u
+  ad=0.81p pd=4.5u as=0p ps=0u
M1221 GND a_626_n285# a_693_n302# Gnd cmosn w=0.9u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1222 VDD a_414_220# S0 w_504_173# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1223 a_359_186# P0 a_323_186# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.81p ps=4.5u
M1224 a_446_67# a_366_79# GND Gnd cmosn w=0.9u l=0.18u
+  ad=0.405p pd=2.7u as=0p ps=0u
M1225 VDD C2 a_653_n135# w_647_n148# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1226 VDD P1 a_203_n209# w_197_n222# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1227 a_57_n598# A3 a_90_n598# Gnd cmosn w=1.8u l=0.18u
+  ad=0.81p pd=4.5u as=0p ps=0u
M1228 a_198_n358# B2 a_162_n358# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.81p ps=4.5u
M1229 VDD A1 a_56_n162# w_50_n175# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1230 a_89_n162# B1 GND Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1231 a_108_98# B0 a_72_98# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.81p ps=4.5u
M1232 a_522_n609# C3 a_486_n609# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.81p ps=4.5u
M1233 a_676_n461# a_587_n446# VDD w_663_n441# cmosp w=1.8u l=0.18u
+  ad=0.81p pd=4.5u as=0p ps=0u
M1234 a_756_n394# P3 GND Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1235 VDD G2 a_723_n394# w_717_n407# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1236 GND A2 a_198_n302# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1237 GND a_162_n302# a_294_n336# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1238 VDD A3 a_72_n518# w_66_n531# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1239 a_162_n104# B1 VDD w_156_n117# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1240 a_330_n175# a_203_n209# a_294_n175# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.81p ps=4.5u
M1241 a_377_n340# P2 VDD w_371_n353# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1242 GND P3 a_431_n587# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1243 C4 a_733_n450# GND Gnd cmosn w=0.9u l=0.18u
+  ad=0.405p pd=2.7u as=0p ps=0u
M1244 a_199_132# a_72_98# a_163_132# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.81p ps=4.5u
M1245 a_562_n169# P2 VDD w_556_n182# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1246 GND a_390_n462# a_733_n450# Gnd cmosn w=0.9u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1247 a_733_n458# a_676_n461# a_733_n466# w_727_n495# cmosp w=9u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1248 a_426_n209# a_294_n231# S1 Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.81p ps=4.5u
M1249 a_409_n332# P1 a_409_n340# Gnd cmosn w=3.6u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1250 a_619_n446# P3 GND Gnd cmosn w=2.7u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1251 a_337_n453# P2 a_337_n461# Gnd cmosn w=2.25u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1252 a_546_n273# P2 VDD w_540_n286# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1253 VDD P2 a_305_n461# w_299_n474# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1254 a_626_n285# a_546_n273# GND Gnd cmosn w=0.9u l=0.18u
+  ad=0.405p pd=2.7u as=0p ps=0u
M1255 GND a_72_n518# a_199_n540# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1256 a_323_186# P0 VDD w_317_173# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1257 a_689_n135# a_562_n169# a_653_n135# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.81p ps=4.5u
M1258 a_239_n209# C1 a_203_n209# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.81p ps=4.5u
M1259 a_57_n598# B3 VDD w_51_n611# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1260 VDD Cin a_414_220# w_408_207# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1261 a_693_n302# a_626_n285# a_693_n310# w_687_n339# cmosp w=7.2u l=0.18u
+  ad=3.24p pd=15.3u as=0p ps=0u
M1262 a_635_n349# a_546_n334# GND Gnd cmosn w=0.9u l=0.18u
+  ad=0.405p pd=2.7u as=0p ps=0u
M1263 a_199_76# B0 a_163_76# Gnd cmosn w=1.8u l=0.18u
+  ad=0p pd=0u as=0.81p ps=4.5u
M1264 VDD a_486_n553# S3 w_576_n600# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1265 a_414_164# P0 VDD w_408_151# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1266 a_404_n97# Cin GND Gnd cmosn w=2.7u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1267 VDD Cin a_377_n340# w_371_n353# cmosp w=1.8u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
.end

