magic
tech scmos
timestamp 1763747745
<< nwell >>
rect -6 16 50 128
<< ntransistor >>
rect 5 0 7 10
rect 13 0 15 10
rect 21 0 23 10
rect 29 0 31 10
rect 37 0 39 10
<< ptransistor >>
rect 5 22 7 122
rect 13 22 15 122
rect 21 22 23 122
rect 29 22 31 122
rect 37 22 39 122
<< ndiffusion >>
rect 4 0 5 10
rect 7 0 8 10
rect 12 0 13 10
rect 15 0 16 10
rect 20 0 21 10
rect 23 0 24 10
rect 28 0 29 10
rect 31 0 32 10
rect 36 0 37 10
rect 39 0 40 10
<< pdiffusion >>
rect 4 22 5 122
rect 7 22 8 122
rect 12 22 13 122
rect 15 22 16 122
rect 20 22 21 122
rect 23 22 24 122
rect 28 22 29 122
rect 31 22 32 122
rect 36 22 37 122
rect 39 22 40 122
<< ndcontact >>
rect 0 0 4 10
rect 8 0 12 10
rect 16 0 20 10
rect 24 0 28 10
rect 32 0 36 10
rect 40 0 44 10
<< pdcontact >>
rect 0 22 4 122
rect 8 22 12 122
rect 16 22 20 122
rect 24 22 28 122
rect 32 22 36 122
rect 40 22 44 122
<< polysilicon >>
rect 5 122 7 131
rect 13 122 15 131
rect 21 122 23 131
rect 29 122 31 131
rect 37 122 39 131
rect 5 10 7 22
rect 13 10 15 22
rect 21 10 23 22
rect 29 10 31 22
rect 37 10 39 22
rect 5 -3 7 0
rect 13 -3 15 0
rect 21 -3 23 0
rect 29 -3 31 0
rect 37 -3 39 0
<< polycontact >>
rect 4 131 8 135
rect 12 131 16 135
rect 20 131 24 135
rect 28 131 32 135
rect 36 131 40 135
<< metal1 >>
rect 4 135 8 139
rect 12 135 16 139
rect 20 135 24 139
rect 28 135 32 139
rect 36 135 40 139
rect -6 125 50 128
rect 0 122 4 125
rect 40 17 44 22
rect 8 16 44 17
rect 8 13 50 16
rect 8 10 12 13
rect 24 10 28 13
rect 40 10 44 13
rect 0 -3 4 0
rect 16 -3 20 0
rect 32 -3 36 0
rect 0 -6 44 -3
rect 47 -9 50 13
<< labels >>
rlabel metal1 -6 125 50 128 1 VDD
rlabel metal1 0 -6 44 -3 1 GND
rlabel metal1 47 -9 50 -6 8 OUT
rlabel metal1 4 135 8 139 5 A
rlabel metal1 12 135 16 139 5 B
rlabel metal1 20 135 24 139 5 C
rlabel metal1 28 135 32 139 5 D
rlabel metal1 36 135 40 139 5 E
<< end >>
