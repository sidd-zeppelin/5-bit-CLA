magic
tech scmos
timestamp 1763728216
<< nwell >>
rect -6 16 18 48
<< ntransistor >>
rect 5 -4 7 6
<< ptransistor >>
rect 5 22 7 42
<< ndiffusion >>
rect 4 -4 5 6
rect 7 -4 8 6
<< pdiffusion >>
rect 4 22 5 42
rect 7 22 8 42
<< ndcontact >>
rect 0 -4 4 6
rect 8 -4 12 6
<< pdcontact >>
rect 0 22 4 42
rect 8 22 12 42
<< polysilicon >>
rect 5 42 7 45
rect 5 6 7 22
rect 5 -7 7 -4
<< polycontact >>
rect 1 9 5 13
<< metal1 >>
rect -6 45 18 48
rect 0 42 4 45
rect 8 13 12 22
rect -6 9 1 13
rect 8 9 18 13
rect 8 6 12 9
rect 0 -7 4 -4
rect 0 -10 12 -7
<< labels >>
rlabel metal1 -6 9 -2 13 3 A
rlabel metal1 14 9 18 13 7 OUT
rlabel metal1 0 -10 12 -7 1 GND
rlabel metal1 -6 45 18 48 5 VDD
<< end >>
