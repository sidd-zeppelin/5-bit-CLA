magic
tech scmos
timestamp 1763745309
<< nwell >>
rect -6 16 42 108
<< ntransistor >>
rect 5 0 7 10
rect 13 0 15 10
rect 21 0 23 10
rect 29 0 31 10
<< ptransistor >>
rect 5 22 7 102
rect 13 22 15 102
rect 21 22 23 102
rect 29 22 31 102
<< ndiffusion >>
rect 4 0 5 10
rect 7 0 8 10
rect 12 0 13 10
rect 15 0 16 10
rect 20 0 21 10
rect 23 0 24 10
rect 28 0 29 10
rect 31 0 32 10
<< pdiffusion >>
rect 4 22 5 102
rect 7 22 8 102
rect 12 22 13 102
rect 15 22 16 102
rect 20 22 21 102
rect 23 22 24 102
rect 28 22 29 102
rect 31 22 32 102
<< ndcontact >>
rect 0 0 4 10
rect 8 0 12 10
rect 16 0 20 10
rect 24 0 28 10
rect 32 0 36 10
<< pdcontact >>
rect 0 22 4 102
rect 8 22 12 102
rect 16 22 20 102
rect 24 22 28 102
rect 32 22 36 102
<< polysilicon >>
rect 5 102 7 111
rect 13 102 15 111
rect 21 102 23 111
rect 29 102 31 111
rect 5 10 7 22
rect 13 10 15 22
rect 21 10 23 22
rect 29 10 31 22
rect 5 -3 7 0
rect 13 -3 15 0
rect 21 -3 23 0
rect 29 -3 31 0
<< polycontact >>
rect 4 111 8 115
rect 12 111 16 115
rect 20 111 24 115
rect 28 111 32 115
<< metal1 >>
rect 4 115 8 119
rect 12 115 16 119
rect 20 115 24 119
rect 28 115 32 119
rect -6 105 42 108
rect 0 102 4 105
rect 32 18 36 22
rect 8 17 36 18
rect 8 14 42 17
rect 8 10 12 14
rect 24 10 28 14
rect 0 -3 4 0
rect 16 -3 20 0
rect 32 -3 36 0
rect 0 -6 36 -3
rect 39 -9 42 14
<< labels >>
rlabel metal1 4 115 8 119 5 A
rlabel metal1 12 115 16 119 5 B
rlabel metal1 20 115 24 119 5 C
rlabel metal1 28 115 32 119 5 D
rlabel metal1 -6 105 42 108 1 VDD
rlabel metal1 0 -6 36 -3 1 GND
rlabel metal1 39 -9 42 -6 8 OUT
<< end >>
