magic
tech scmos
timestamp 1764587577
<< nwell >>
rect 6 -55 28 9
<< ntransistor >>
rect 36 -4 66 -2
rect 36 -12 66 -10
rect 36 -20 66 -18
rect 36 -28 66 -26
rect 36 -36 66 -34
rect 36 -44 66 -42
<< ptransistor >>
rect 12 -4 22 -2
rect 12 -12 22 -10
rect 12 -20 22 -18
rect 12 -28 22 -26
rect 12 -36 22 -34
rect 12 -44 22 -42
<< ndiffusion >>
rect 36 -2 66 -1
rect 36 -5 66 -4
rect 36 -10 66 -9
rect 36 -13 66 -12
rect 36 -18 66 -17
rect 36 -21 66 -20
rect 36 -26 66 -25
rect 36 -29 66 -28
rect 36 -34 66 -33
rect 36 -37 66 -36
rect 36 -42 66 -41
rect 36 -45 66 -44
<< pdiffusion >>
rect 12 -2 22 -1
rect 12 -5 22 -4
rect 12 -10 22 -9
rect 12 -13 22 -12
rect 12 -18 22 -17
rect 12 -21 22 -20
rect 12 -26 22 -25
rect 12 -29 22 -28
rect 12 -34 22 -33
rect 12 -37 22 -36
rect 12 -42 22 -41
rect 12 -45 22 -44
<< ndcontact >>
rect 36 -1 66 3
rect 36 -9 66 -5
rect 36 -17 66 -13
rect 36 -25 66 -21
rect 36 -33 66 -29
rect 36 -41 66 -37
rect 36 -49 66 -45
<< pdcontact >>
rect 12 -1 22 3
rect 12 -9 22 -5
rect 12 -17 22 -13
rect 12 -25 22 -21
rect 12 -33 22 -29
rect 12 -41 22 -37
rect 12 -49 22 -45
<< polysilicon >>
rect 2 -4 12 -2
rect 22 -4 36 -2
rect 66 -4 69 -2
rect 2 -12 12 -10
rect 22 -12 36 -10
rect 66 -12 69 -10
rect 2 -20 12 -18
rect 22 -20 36 -18
rect 66 -20 69 -18
rect 2 -28 12 -26
rect 22 -28 36 -26
rect 66 -28 69 -26
rect 2 -36 12 -34
rect 22 -36 36 -34
rect 66 -36 69 -34
rect 2 -44 12 -42
rect 22 -44 36 -42
rect 66 -44 69 -42
<< polycontact >>
rect -2 -5 2 -1
rect -2 -13 2 -9
rect -2 -21 2 -17
rect -2 -29 2 -25
rect -2 -37 2 -33
rect -2 -45 2 -41
<< metal1 >>
rect 5 3 9 9
rect 28 6 77 10
rect 28 3 32 6
rect 5 -1 12 3
rect 28 -1 36 3
rect -6 -5 -2 -1
rect -6 -13 -2 -9
rect 5 -13 9 -1
rect 28 -5 32 -1
rect 22 -9 32 -5
rect 5 -17 12 -13
rect -6 -21 -2 -17
rect -6 -29 -2 -25
rect 5 -29 9 -17
rect 28 -21 32 -9
rect 22 -25 32 -21
rect 5 -33 12 -29
rect -6 -37 -2 -33
rect -6 -45 -2 -41
rect 5 -45 9 -33
rect 28 -37 32 -25
rect 22 -41 32 -37
rect 69 -45 73 3
rect 5 -49 12 -45
rect 66 -49 73 -45
rect 5 -55 9 -49
<< labels >>
rlabel metal1 69 -49 73 3 7 GND
rlabel metal1 5 -55 9 9 3 VDD
rlabel metal1 -6 -45 -2 -41 3 A
rlabel metal1 -6 -37 -2 -33 3 B
rlabel metal1 -6 -29 -2 -25 3 C
rlabel metal1 -6 -21 -2 -17 3 D
rlabel metal1 -6 -13 -2 -9 3 E
rlabel metal1 -6 -5 -2 -1 3 F
rlabel metal1 73 6 77 10 6 OUT
<< end >>
