magic
tech scmos
timestamp 1763641429
<< nwell >>
rect 105 34 137 66
rect 14 0 46 32
rect 105 -22 137 10
rect 201 0 233 32
<< ntransistor >>
rect 147 53 167 55
rect 147 45 167 47
rect 56 19 76 21
rect 243 19 263 21
rect 56 11 76 13
rect 243 11 263 13
rect 147 -3 167 -1
rect 147 -11 167 -9
<< ptransistor >>
rect 111 53 131 55
rect 111 45 131 47
rect 20 19 40 21
rect 207 19 227 21
rect 20 11 40 13
rect 207 11 227 13
rect 111 -3 131 -1
rect 111 -11 131 -9
<< ndiffusion >>
rect 147 55 167 56
rect 147 52 167 53
rect 147 47 167 48
rect 147 44 167 45
rect 56 21 76 22
rect 56 18 76 19
rect 243 21 263 22
rect 56 13 76 14
rect 56 10 76 11
rect 243 18 263 19
rect 243 13 263 14
rect 243 10 263 11
rect 147 -1 167 0
rect 147 -4 167 -3
rect 147 -9 167 -8
rect 147 -12 167 -11
<< pdiffusion >>
rect 111 55 131 56
rect 111 52 131 53
rect 111 47 131 48
rect 111 44 131 45
rect 20 21 40 22
rect 20 18 40 19
rect 20 13 40 14
rect 207 21 227 22
rect 207 18 227 19
rect 20 10 40 11
rect 207 13 227 14
rect 207 10 227 11
rect 111 -1 131 0
rect 111 -4 131 -3
rect 111 -9 131 -8
rect 111 -12 131 -11
<< ndcontact >>
rect 147 56 167 60
rect 147 48 167 52
rect 147 40 167 44
rect 56 22 76 26
rect 243 22 263 26
rect 56 14 76 18
rect 243 14 263 18
rect 56 6 76 10
rect 243 6 263 10
rect 147 0 167 4
rect 147 -8 167 -4
rect 147 -16 167 -12
<< pdcontact >>
rect 111 56 131 60
rect 111 48 131 52
rect 111 40 131 44
rect 20 22 40 26
rect 207 22 227 26
rect 20 14 40 18
rect 207 14 227 18
rect 20 6 40 10
rect 207 6 227 10
rect 111 0 131 4
rect 111 -8 131 -4
rect 111 -16 131 -12
<< polysilicon >>
rect 99 53 111 55
rect 131 53 147 55
rect 167 53 170 55
rect 99 45 111 47
rect 131 45 147 47
rect 167 45 170 47
rect 8 19 20 21
rect 40 19 56 21
rect 76 19 79 21
rect 195 19 207 21
rect 227 19 243 21
rect 263 19 266 21
rect 8 11 20 13
rect 40 11 56 13
rect 76 11 79 13
rect 195 11 207 13
rect 227 11 243 13
rect 263 11 266 13
rect 99 -3 111 -1
rect 131 -3 147 -1
rect 167 -3 170 -1
rect 99 -11 111 -9
rect 131 -11 147 -9
rect 167 -11 170 -9
<< polycontact >>
rect 95 52 99 56
rect 95 44 99 48
rect 4 18 8 22
rect 4 10 8 14
rect 191 18 195 22
rect 191 10 195 14
rect 95 -4 99 0
rect 95 -12 99 -8
<< metal1 >>
rect -12 74 201 78
rect 139 63 182 67
rect 102 56 111 60
rect 0 52 95 56
rect 0 22 4 52
rect 91 33 95 48
rect 102 44 105 56
rect 139 52 143 63
rect 167 56 170 60
rect 131 48 143 52
rect 139 44 143 48
rect 48 29 95 33
rect 11 22 20 26
rect -12 18 4 22
rect -12 10 4 14
rect 11 10 14 22
rect 48 18 52 29
rect 76 22 80 26
rect 40 14 52 18
rect 48 10 52 14
rect 0 -8 4 10
rect 11 6 20 10
rect 48 6 56 10
rect 91 -4 95 29
rect 102 40 111 44
rect 139 40 147 44
rect 102 31 106 40
rect 102 27 151 31
rect 102 4 106 27
rect 178 22 182 63
rect 197 31 201 74
rect 235 30 285 34
rect 198 22 207 26
rect 178 18 191 22
rect 178 11 191 14
rect 139 10 191 11
rect 198 10 201 22
rect 235 18 239 30
rect 263 22 267 26
rect 227 14 239 18
rect 235 10 239 14
rect 139 7 182 10
rect 102 0 111 4
rect 0 -12 95 -8
rect 102 -12 105 0
rect 139 -4 143 7
rect 198 6 207 10
rect 235 6 243 10
rect 167 0 177 4
rect 131 -8 143 -4
rect 139 -12 143 -8
rect 102 -16 111 -12
rect 139 -16 147 -12
rect 173 -19 177 0
rect 267 -19 271 22
rect -12 -23 271 -19
<< m2contact >>
rect 10 69 15 74
rect 170 55 175 60
rect 10 26 15 31
rect 80 21 85 26
rect 151 27 156 32
rect 196 26 201 31
rect 267 22 272 27
<< metal2 >>
rect 11 31 14 69
rect 172 48 175 55
rect 172 45 271 48
rect 172 39 175 45
rect 144 36 175 39
rect 144 25 147 36
rect 156 28 196 31
rect 268 27 271 45
rect 85 22 147 25
<< labels >>
rlabel metal1 281 30 285 34 7 OUT
rlabel metal1 -12 18 -8 22 3 A
rlabel metal1 -12 10 -8 14 3 B
rlabel metal1 -12 74 -8 78 4 VDD
rlabel metal1 -12 -23 -8 -19 2 GND
<< end >>
