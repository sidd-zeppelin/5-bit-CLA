magic
tech scmos
timestamp 1764717201
<< nwell >>
rect 11 0 63 32
rect 94 22 118 54
<< polysilicon >>
rect 105 48 107 51
rect 8 19 17 21
rect 57 19 69 21
rect 79 19 82 21
rect 8 11 17 13
rect 57 11 69 13
rect 79 11 82 13
rect 105 12 107 28
rect 105 -1 107 2
<< ndiffusion >>
rect 69 21 79 22
rect 69 18 79 19
rect 69 13 79 14
rect 69 10 79 11
rect 104 2 105 12
rect 107 2 108 12
<< pdiffusion >>
rect 104 28 105 48
rect 107 28 108 48
rect 17 21 57 22
rect 17 18 57 19
rect 17 13 57 14
rect 17 10 57 11
<< metal1 >>
rect 0 51 118 54
rect 0 18 4 22
rect 0 10 4 14
rect 11 10 14 51
rect 100 48 104 51
rect 63 29 91 32
rect 63 26 66 29
rect 57 22 66 26
rect 79 22 85 26
rect 63 18 66 22
rect 63 14 69 18
rect 82 10 85 22
rect 88 19 91 29
rect 108 19 112 28
rect 88 15 101 19
rect 108 15 118 19
rect 108 12 112 15
rect 11 6 17 10
rect 79 6 85 10
rect 82 -1 85 6
rect 100 -1 104 2
rect 0 -4 112 -1
<< ntransistor >>
rect 69 19 79 21
rect 69 11 79 13
rect 105 2 107 12
<< ptransistor >>
rect 105 28 107 48
rect 17 19 57 21
rect 17 11 57 13
<< polycontact >>
rect 4 18 8 22
rect 4 10 8 14
rect 101 15 105 19
<< ndcontact >>
rect 69 22 79 26
rect 69 14 79 18
rect 69 6 79 10
rect 100 2 104 12
rect 108 2 112 12
<< pdcontact >>
rect 100 28 104 48
rect 108 28 112 48
rect 17 22 57 26
rect 17 14 57 18
rect 17 6 57 10
<< labels >>
rlabel metal1 0 10 4 14 3 A
rlabel metal1 0 18 4 22 3 B
rlabel metal1 114 15 118 19 7 OUT
rlabel metal1 0 51 3 54 4 VDD
rlabel metal1 0 -4 3 -1 2 GND
<< end >>
