* NGSPICE file created from NAND6.ext - technology: scmos

.global Vdd Gnd 


* Top level circuit NAND6

M1000 a_39_n44# E a_31_n44# Gnd cmosn w=2.7u l=0.18u
+  ad=1.458p pd=6.48u as=1.458p ps=6.48u
M1001 VDD D OUT w_n6_n6# cmosp w=0.9u l=0.18u
+  ad=1.782p pd=11.16u as=1.458p ps=8.64u
M1002 VDD B OUT w_n6_n6# cmosp w=0.9u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1003 OUT F a_39_n44# Gnd cmosn w=2.7u l=0.18u
+  ad=1.215p pd=6.3u as=0p ps=0u
M1004 OUT A VDD w_n6_n6# cmosp w=0.9u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1005 OUT E VDD w_n6_n6# cmosp w=0.9u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1006 OUT C VDD w_n6_n6# cmosp w=0.9u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1007 VDD F OUT w_n6_n6# cmosp w=0.9u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1008 a_15_n44# B a_7_n44# Gnd cmosn w=2.7u l=0.18u
+  ad=1.458p pd=6.48u as=1.458p ps=6.48u
M1009 a_7_n44# A GND Gnd cmosn w=2.7u l=0.18u
+  ad=0p pd=0u as=1.215p ps=6.3u
M1010 a_31_n44# D a_23_n44# Gnd cmosn w=2.7u l=0.18u
+  ad=0p pd=0u as=1.458p ps=6.48u
M1011 a_23_n44# C a_15_n44# Gnd cmosn w=2.7u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
.end

