* NGSPICE file created from AND6.ext - technology: scmos

.global Vdd Gnd 


* Top level circuit AND6

M1000 VDD D a_18_13# w_11_0# cmosp w=0.9u l=0.18u
+  ad=2.592p pd=15.66u as=1.458p ps=8.64u
M1001 a_18_13# F a_42_45# Gnd cmosn w=2.7u l=0.18u
+  ad=1.215p pd=6.3u as=1.458p ps=6.48u
M1002 a_42_29# C a_42_21# Gnd cmosn w=2.7u l=0.18u
+  ad=1.458p pd=6.48u as=1.458p ps=6.48u
M1003 a_18_13# E VDD w_11_0# cmosp w=0.9u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1004 a_42_13# A GND Gnd cmosn w=2.7u l=0.18u
+  ad=1.458p pd=6.48u as=1.62p ps=9u
M1005 VDD B a_18_13# w_11_0# cmosp w=0.9u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1006 OUT a_18_13# GND Gnd cmosn w=0.9u l=0.18u
+  ad=0.405p pd=2.7u as=0p ps=0u
M1007 a_42_37# D a_42_29# Gnd cmosn w=2.7u l=0.18u
+  ad=1.458p pd=6.48u as=0p ps=0u
M1008 VDD F a_18_13# w_11_0# cmosp w=0.9u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1009 OUT a_18_13# VDD w_93_33# cmosp w=1.8u l=0.18u
+  ad=0.81p pd=4.5u as=0p ps=0u
M1010 a_18_13# C VDD w_11_0# cmosp w=0.9u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1011 a_42_45# E a_42_37# Gnd cmosn w=2.7u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1012 a_42_21# B a_42_13# Gnd cmosn w=2.7u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
M1013 a_18_13# A VDD w_11_0# cmosp w=0.9u l=0.18u
+  ad=0p pd=0u as=0p ps=0u
.end

