magic
tech scmos
timestamp 1763602483
<< nwell >>
rect -28 -14 4 18
rect 78 4 110 36
rect 299 -14 331 18
rect 405 4 437 36
rect -124 -46 -100 -14
rect -73 -46 -49 -14
rect -28 -61 4 -29
rect 78 -61 110 -29
rect 204 -46 228 -14
rect 254 -46 278 -14
rect 299 -61 331 -29
rect 405 -61 437 -29
<< ntransistor >>
rect 120 23 140 25
rect 447 23 467 25
rect 120 15 140 17
rect 447 15 467 17
rect 14 5 34 7
rect 341 5 361 7
rect 14 -3 34 -1
rect 341 -3 361 -1
rect 14 -42 34 -40
rect 120 -42 140 -40
rect 14 -50 34 -48
rect -113 -64 -111 -54
rect -62 -64 -60 -54
rect 120 -50 140 -48
rect 341 -42 361 -40
rect 447 -42 467 -40
rect 341 -50 361 -48
rect 215 -64 217 -54
rect 265 -64 267 -54
rect 447 -50 467 -48
<< ptransistor >>
rect 84 23 104 25
rect 411 23 431 25
rect 84 15 104 17
rect 411 15 431 17
rect -22 5 -2 7
rect 305 5 325 7
rect -22 -3 -2 -1
rect 305 -3 325 -1
rect -113 -40 -111 -20
rect -62 -40 -60 -20
rect -22 -42 -2 -40
rect 215 -40 217 -20
rect 265 -40 267 -20
rect 84 -42 104 -40
rect -22 -50 -2 -48
rect 84 -50 104 -48
rect 305 -42 325 -40
rect 411 -42 431 -40
rect 305 -50 325 -48
rect 411 -50 431 -48
<< ndiffusion >>
rect 120 25 140 26
rect 120 22 140 23
rect 447 25 467 26
rect 120 17 140 18
rect 120 14 140 15
rect 447 22 467 23
rect 447 17 467 18
rect 14 7 34 8
rect 14 4 34 5
rect 447 14 467 15
rect 341 7 361 8
rect 14 -1 34 0
rect 14 -4 34 -3
rect 341 4 361 5
rect 341 -1 361 0
rect 341 -4 361 -3
rect 14 -40 34 -39
rect 14 -43 34 -42
rect 120 -40 140 -39
rect 14 -48 34 -47
rect -114 -64 -113 -54
rect -111 -64 -110 -54
rect -63 -64 -62 -54
rect -60 -64 -59 -54
rect 14 -51 34 -50
rect 120 -43 140 -42
rect 120 -48 140 -47
rect 120 -51 140 -50
rect 341 -40 361 -39
rect 341 -43 361 -42
rect 447 -40 467 -39
rect 341 -48 361 -47
rect 214 -64 215 -54
rect 217 -64 218 -54
rect 264 -64 265 -54
rect 267 -64 268 -54
rect 341 -51 361 -50
rect 447 -43 467 -42
rect 447 -48 467 -47
rect 447 -51 467 -50
<< pdiffusion >>
rect 84 25 104 26
rect 84 22 104 23
rect 84 17 104 18
rect 411 25 431 26
rect 411 22 431 23
rect 84 14 104 15
rect -22 7 -2 8
rect 411 17 431 18
rect 411 14 431 15
rect -22 4 -2 5
rect -22 -1 -2 0
rect 305 7 325 8
rect 305 4 325 5
rect -22 -4 -2 -3
rect 305 -1 325 0
rect 305 -4 325 -3
rect -114 -40 -113 -20
rect -111 -40 -110 -20
rect -63 -40 -62 -20
rect -60 -40 -59 -20
rect -22 -40 -2 -39
rect -22 -43 -2 -42
rect -22 -48 -2 -47
rect 84 -40 104 -39
rect 214 -40 215 -20
rect 217 -40 218 -20
rect 264 -40 265 -20
rect 267 -40 268 -20
rect 84 -43 104 -42
rect -22 -51 -2 -50
rect 84 -48 104 -47
rect 84 -51 104 -50
rect 305 -40 325 -39
rect 305 -43 325 -42
rect 305 -48 325 -47
rect 411 -40 431 -39
rect 411 -43 431 -42
rect 305 -51 325 -50
rect 411 -48 431 -47
rect 411 -51 431 -50
<< ndcontact >>
rect 120 26 140 30
rect 447 26 467 30
rect 120 18 140 22
rect 14 8 34 12
rect 447 18 467 22
rect 120 10 140 14
rect 341 8 361 12
rect 447 10 467 14
rect 14 0 34 4
rect 341 0 361 4
rect 14 -8 34 -4
rect 341 -8 361 -4
rect 14 -39 34 -35
rect 120 -39 140 -35
rect 14 -47 34 -43
rect -118 -64 -114 -54
rect -110 -64 -106 -54
rect -67 -64 -63 -54
rect -59 -64 -55 -54
rect 120 -47 140 -43
rect 14 -55 34 -51
rect 120 -55 140 -51
rect 341 -39 361 -35
rect 447 -39 467 -35
rect 341 -47 361 -43
rect 210 -64 214 -54
rect 218 -64 222 -54
rect 260 -64 264 -54
rect 268 -64 272 -54
rect 447 -47 467 -43
rect 341 -55 361 -51
rect 447 -55 467 -51
<< pdcontact >>
rect 84 26 104 30
rect 411 26 431 30
rect 84 18 104 22
rect 411 18 431 22
rect -22 8 -2 12
rect 84 10 104 14
rect 305 8 325 12
rect -22 0 -2 4
rect 411 10 431 14
rect 305 0 325 4
rect -22 -8 -2 -4
rect 305 -8 325 -4
rect -118 -40 -114 -20
rect -110 -40 -106 -20
rect -67 -40 -63 -20
rect -59 -40 -55 -20
rect -22 -39 -2 -35
rect 84 -39 104 -35
rect -22 -47 -2 -43
rect 210 -40 214 -20
rect 218 -40 222 -20
rect 260 -40 264 -20
rect 268 -40 272 -20
rect 305 -39 325 -35
rect 84 -47 104 -43
rect -22 -55 -2 -51
rect 84 -55 104 -51
rect 411 -39 431 -35
rect 305 -47 325 -43
rect 411 -47 431 -43
rect 305 -55 325 -51
rect 411 -55 431 -51
<< polysilicon >>
rect 72 23 84 25
rect 104 23 120 25
rect 140 23 143 25
rect 399 23 411 25
rect 431 23 447 25
rect 467 23 470 25
rect 72 15 84 17
rect 104 15 120 17
rect 140 15 143 17
rect 399 15 411 17
rect 431 15 447 17
rect 467 15 470 17
rect -34 5 -22 7
rect -2 5 14 7
rect 34 5 37 7
rect 293 5 305 7
rect 325 5 341 7
rect 361 5 364 7
rect -34 -3 -22 -1
rect -2 -3 14 -1
rect 34 -3 37 -1
rect 293 -3 305 -1
rect 325 -3 341 -1
rect 361 -3 364 -1
rect -113 -20 -111 -17
rect -62 -20 -60 -17
rect 215 -20 217 -17
rect 265 -20 267 -17
rect -113 -54 -111 -40
rect -62 -54 -60 -40
rect -34 -42 -22 -40
rect -2 -42 14 -40
rect 34 -42 37 -40
rect 72 -42 84 -40
rect 104 -42 120 -40
rect 140 -42 143 -40
rect -34 -50 -22 -48
rect -2 -50 14 -48
rect 34 -50 37 -48
rect 72 -50 84 -48
rect 104 -50 120 -48
rect 140 -50 143 -48
rect 215 -54 217 -40
rect 265 -54 267 -40
rect 293 -42 305 -40
rect 325 -42 341 -40
rect 361 -42 364 -40
rect 399 -42 411 -40
rect 431 -42 447 -40
rect 467 -42 470 -40
rect 293 -50 305 -48
rect 325 -50 341 -48
rect 361 -50 364 -48
rect 399 -50 411 -48
rect 431 -50 447 -48
rect 467 -50 470 -48
rect -113 -67 -111 -64
rect -62 -67 -60 -64
rect 215 -67 217 -64
rect 265 -67 267 -64
<< polycontact >>
rect 68 22 72 26
rect 68 14 72 18
rect 395 22 399 26
rect -38 4 -34 8
rect 395 14 399 18
rect -38 -4 -34 0
rect 289 4 293 8
rect 289 -4 293 0
rect -117 -51 -113 -47
rect -66 -51 -62 -47
rect -38 -43 -34 -39
rect -38 -51 -34 -47
rect 68 -43 72 -39
rect 68 -51 72 -47
rect 211 -51 215 -47
rect 261 -51 265 -47
rect 289 -43 293 -39
rect 289 -51 293 -47
rect 395 -43 399 -39
rect 395 -51 399 -47
<< metal1 >>
rect 26 47 300 50
rect 26 44 29 47
rect 296 44 300 47
rect -124 41 78 44
rect -31 12 -28 41
rect 75 30 78 41
rect 296 41 405 44
rect 112 36 248 40
rect 75 26 84 30
rect 6 22 68 26
rect -31 8 -22 12
rect -139 4 -38 8
rect -124 -14 -104 -10
rect -118 -20 -114 -14
rect -110 -47 -106 -40
rect -93 -47 -90 -5
rect -139 -51 -117 -47
rect -110 -51 -90 -47
rect -83 -47 -79 4
rect -68 -14 -54 -10
rect -67 -20 -63 -14
rect -59 -47 -55 -40
rect -42 -43 -38 0
rect -31 -4 -28 8
rect 6 4 10 22
rect 40 12 43 18
rect 34 8 43 12
rect -2 0 10 4
rect 6 -4 10 0
rect -31 -8 -22 -4
rect 6 -8 14 -4
rect -31 -11 -28 -8
rect 40 -10 43 8
rect 75 14 78 26
rect 112 22 116 36
rect 140 26 142 30
rect 104 18 116 22
rect 112 14 116 18
rect 68 7 71 14
rect 75 10 84 14
rect 112 10 120 14
rect 75 4 78 10
rect 150 -1 154 36
rect 68 -5 154 -1
rect 6 -25 52 -21
rect -31 -35 -28 -32
rect -31 -39 -22 -35
rect -83 -51 -66 -47
rect -59 -51 -38 -47
rect -31 -51 -28 -39
rect 6 -43 10 -25
rect 40 -35 43 -33
rect 34 -39 43 -35
rect -2 -47 10 -43
rect 6 -51 10 -47
rect -110 -54 -106 -51
rect -59 -54 -55 -51
rect -31 -55 -22 -51
rect 6 -55 14 -51
rect -31 -61 -28 -55
rect -118 -70 -114 -64
rect -67 -70 -63 -64
rect 40 -70 43 -39
rect 48 -47 52 -25
rect 68 -39 72 -5
rect 75 -35 78 -29
rect 75 -39 84 -35
rect 48 -51 68 -47
rect 75 -51 78 -39
rect 112 -43 116 -13
rect 160 -35 163 26
rect 244 8 248 36
rect 296 12 299 41
rect 402 30 405 41
rect 439 36 513 40
rect 402 26 411 30
rect 333 22 395 26
rect 296 8 305 12
rect 244 4 289 8
rect 204 -14 228 -10
rect 140 -39 163 -35
rect 104 -47 116 -43
rect 112 -51 116 -47
rect 75 -55 84 -51
rect 112 -55 120 -51
rect 75 -61 78 -55
rect 160 -70 163 -39
rect 210 -20 214 -14
rect 218 -47 222 -40
rect 234 -47 239 -5
rect 199 -51 211 -47
rect 218 -51 239 -47
rect 244 -47 248 4
rect 259 -14 273 -10
rect 260 -20 264 -14
rect 268 -47 272 -40
rect 285 -43 289 0
rect 296 -4 299 8
rect 333 4 337 22
rect 367 12 370 18
rect 361 8 370 12
rect 325 0 337 4
rect 333 -4 337 0
rect 296 -8 305 -4
rect 333 -8 341 -4
rect 296 -11 299 -8
rect 367 -10 370 8
rect 402 14 405 26
rect 439 22 443 36
rect 467 26 469 30
rect 431 18 443 22
rect 439 14 443 18
rect 395 7 398 14
rect 402 10 411 14
rect 439 10 447 14
rect 402 4 405 10
rect 477 -1 481 36
rect 395 -5 481 -1
rect 333 -25 379 -21
rect 296 -35 299 -32
rect 296 -39 305 -35
rect 244 -51 261 -47
rect 268 -51 289 -47
rect 296 -51 299 -39
rect 333 -43 337 -25
rect 367 -35 370 -33
rect 361 -39 370 -35
rect 325 -47 337 -43
rect 333 -51 337 -47
rect 218 -54 222 -51
rect 268 -54 272 -51
rect 296 -55 305 -51
rect 333 -55 341 -51
rect 296 -61 299 -55
rect 210 -70 214 -64
rect 260 -70 264 -64
rect 367 -70 370 -39
rect 375 -47 379 -25
rect 395 -39 399 -5
rect 402 -35 405 -29
rect 402 -39 411 -35
rect 375 -51 395 -47
rect 402 -51 405 -39
rect 439 -43 443 -13
rect 487 -35 490 26
rect 467 -39 490 -35
rect 431 -47 443 -43
rect 439 -51 443 -47
rect 402 -55 411 -51
rect 439 -55 447 -51
rect 402 -61 405 -55
rect 487 -70 490 -39
rect -118 -73 490 -70
<< m2contact >>
rect 58 36 63 41
rect -94 -5 -89 0
rect -104 -14 -99 -9
rect -47 -5 -42 0
rect -73 -14 -68 -9
rect -54 -14 -49 -9
rect 142 26 147 31
rect 66 2 71 7
rect 111 2 117 7
rect 159 26 164 31
rect -33 -16 -28 -11
rect 39 -15 44 -10
rect -33 -32 -28 -27
rect 40 -33 45 -28
rect 111 -13 117 -8
rect 75 -29 80 -24
rect 291 18 296 24
rect 385 36 390 41
rect 234 -5 239 0
rect 216 -10 221 -5
rect 194 -52 199 -47
rect 280 -5 285 0
rect 254 -14 259 -9
rect 273 -14 278 -9
rect 469 26 474 31
rect 393 2 398 7
rect 438 2 444 7
rect 486 26 491 31
rect 294 -16 299 -11
rect 366 -15 371 -10
rect 294 -32 299 -27
rect 367 -33 372 -28
rect 438 -13 444 -8
rect 402 -29 407 -24
<< metal2 >>
rect -59 51 198 54
rect -59 -1 -56 51
rect -89 -4 -47 -1
rect -99 -13 -73 -10
rect -49 -14 -33 -11
rect -33 -27 -28 -16
rect 40 -28 43 -15
rect 59 -25 62 36
rect 147 27 159 30
rect 71 2 111 5
rect 112 -8 116 2
rect 59 -28 75 -25
rect 195 -47 198 51
rect 217 19 291 22
rect 217 -5 220 19
rect 239 -4 280 -1
rect 278 -14 294 -11
rect 295 -27 298 -16
rect 367 -28 370 -15
rect 386 -25 389 36
rect 474 27 486 30
rect 398 2 438 5
rect 439 -8 443 2
rect 386 -28 402 -25
<< labels >>
rlabel metal1 -139 4 -135 8 3 D_in
rlabel metal1 -139 -51 -135 -47 3 CLK
rlabel metal1 -118 -73 -114 -70 1 GND
rlabel metal1 -124 41 -121 44 1 VDD
rlabel metal1 508 36 513 40 7 Q
<< end >>
